.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.param width_N={10*LAMBDA}
.param width_P={20*LAMBDA}
.global gnd vdd

Vdd vdd gnd 'SUPPLY'
vd10 a1in 0 pulse 1.8 0 0ns 100ps 100ps 9.8ns 29.8ns
vd_bar10 a1in_inv 0 pulse 0 1.8 0ns 100ps 100ps 9.8ns 29.8ns
vd11 b1in_inv 0 pulse 1.8 0 0ns 100ps 100ps 9.8ns 29.8ns
vd_bar11 b1in 0 pulse 0 1.8 0ns 100ps 100ps 9.8ns 29.8ns
vclk clk 0 pulse 1.8 0 0ns 100ps 100ps 10ns 20ns




* INVERTER
.subckt inv x y vdd gnd
M1 y x gnd gnd CMOSN W={width_N} L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA}
PD={10*LAMBDA+2*width_N}
M2 y x vdd vdd CMOSP W={width_P} L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA}
PD={10*LAMBDA+2*width_P}
.ends inv
* NAND, Note that this is only used for Dlatch and flipflop
.subckt nand x1 x2 y vdd gnd
M1 y x2 vdd vdd CMOSP W={width_P} L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA}
PD={10*LAMBDA+2*width_P}
M2 y x1 vdd vdd CMOSP W={width_P} L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA}
PD={10*LAMBDA+2*width_P}
M3 y x1 xbtw xbtw CMOSN W={2*width_N} L={2*LAMBDA}
+ AS={5*2*width_N*LAMBDA} PS={10*LAMBDA+2*2*width_N} AD={5*2*width_N*LAMBDA}
PD={10*LAMBDA+2*2*width_N}
M4 xbtw x2 gnd gnd CMOSN W={2*width_N} L={2*LAMBDA}
+ AS={5*2*width_N*LAMBDA} PS={10*LAMBDA+2*2*width_N} AD={5*2*width_N*LAMBDA}
PD={10*LAMBDA+2*2*width_N}
.ends nand
* Dlatch, Note that this is only used to make the flipflop
.subckt dlatch enable d d_inv q q_inv vdd gnd
xx1 enable d s vdd gnd nand
xx2 enable d_inv r vdd gnd nand
xx3 s q_inv q vdd gnd nand
xx4 r q q_inv vdd gnd nand
.ends dlatch
*Dflipflop, used twice in the final circuit
.subckt dflipflop clk d d_inv q q_inv vdd gnd
xxx3 clk clk_inv vdd gnd inv
xxx1 clk_inv d d_inv xbtw xbtw_inv vdd gnd dlatch
xxx2 clk xbtw xbtw_inv q q_inv vdd gnd dlatch
.ends dflipflop


x1 clk a1in a1in_inv a1 a1_inv vdd gnd dflipflop
x2 clk b1in b1in_inv b1 b1_inv vdd gnd dflipflop

.tran 2ps 40n
.control
set hcopypscolor = 1
set color0=white
set color1=black
run
set curplottitle= "Abhayram A Nair-2019102017"
plot v(a1in) v(a1)+2 v(clk)+4
set curplottitle= "Abhayram A Nair-2019102017"
plot v(b1in) v(b1)+2 v(clk)+4
.endc