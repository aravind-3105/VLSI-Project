* SPICE3 file created from xorlabel.ext - technology: scmos

.option scale=0.09u

M1000 a_80_n16# x2 vdd inv_1/w_n16_11# pfet w=20 l=2
+  ad=100 pd=50 as=440 ps=192
M1001 a_80_n16# x2 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=300 ps=160
M1002 a_72_n5# x1 vdd inv_0/w_n16_11# pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1003 a_72_n5# x1 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1004 vdd x1 a_53_26# w_47_20# pfet w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M1005 a_53_26# x2 vdd w_47_20# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 y a_72_n5# a_53_26# w_47_20# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1007 a_53_26# a_80_n16# y w_47_20# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1008 a_60_n47# x1 gnd Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1009 y x2 a_60_n47# Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1010 a_76_n47# a_72_n5# y Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1011 gnd a_80_n16# a_76_n47# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
C0 x2 x1 1.7fF
C1 w_47_20# gnd! 2.5fF
C2 vdd gnd! 1.3fF
C3 gnd gnd! 1.6fF
