* SPICE3 file created from 3AND.ext - technology: scmos

.option scale=0.09u

M1000 out C vdd w_0_0# pfet w=20 l=2
+  ad=220 pd=102 as=220 ps=102
M1001 vdd B out w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 out A vdd w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 a_13_n61# C gnd Gnd nfet w=30 l=2
+  ad=180 pd=72 as=150 ps=70
M1004 a_21_n61# B a_13_n61# Gnd nfet w=30 l=2
+  ad=180 pd=72 as=0 ps=0
M1005 out A a_21_n61# Gnd nfet w=30 l=2
+  ad=210 pd=74 as=0 ps=0
C0 w_0_0# gnd! 1.5fF
