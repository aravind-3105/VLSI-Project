.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.param width_N={20*LAMBDA}
.param width_P={40*LAMBDA}
.global gnd vdd

Vdd	vdd	gnd	'SUPPLY'
vd1 a 0 pulse 1.8 0 0ns 100ps 100ps 10ns 60ns
vd2 b 0 pulse 0 1.8 0ns 100ps 100ps 20ns 60ns






.subckt and_subckt a b y vdd gnd
* Layer-1
M1      nand       b       vdd     vdd  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

M2      nand       a       vdd     vdd  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}


M3      nand       a       J     J  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

M4      J         b      gnd gnd   CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}


M5      y       nand       vdd     vdd  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

M6      y       nand       gnd     gnd  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
.ends and_subckt

x1 a b y vdd gnd and_subckt

.tran 1n 60n


.control
set hcopypscolor = 1
set color0=white
set color1=black

run
plot v(a)
plot v(b)
plot v(y)
set curplottitle= "Aravind Narayanan-2019102014"
.endc