* SPICE3 file created from 3AND.ext - technology: scmos
.option scale=0.09u
.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.global gnd vdd

Vdd	vdd	gnd	'SUPPLY'
vdA     A     0 pulse 1.8 0 0ns 100ps 100ps 5ns  30ns
vdB     B     0 pulse 1.8 0 30ns 100ps 100ps 10ns  30ns
vdC     C     0 pulse 1.8 0 30ns 100ps 100ps 20ns  40ns

M1000 a_14_3# C vdd w_1_n3# CMOSP w=60 l=2
+  ad=360 pd=132 as=300 ps=130
M1001 a_22_3# B a_14_3# w_1_n3# CMOSP w=60 l=2
+  ad=360 pd=132 as=0 ps=0
M1002 out A a_22_3# w_1_n3# CMOSP w=60 l=2
+  ad=420 pd=134 as=0 ps=0
M1003 out C gnd gnd CMOSN w=10 l=2
+  ad=130 pd=66 as=110 ps=62
M1004 gnd B out gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 out A gnd gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
C0 w_1_n3# gnd 3.3fF





.tran 1n 60n
.control
set hcopypscolor = 1
set color0=white
set color1=black

run
plot v(A) v(B)+2 v(C)+4 v(out)+8
set curplottitle= "Aravind Narayanan-2019102014"
.endc