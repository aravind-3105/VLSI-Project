* SPICE3 file created from 4AND.ext - technology: scmos

.option scale=0.09u

M1000 out D vdd w_0_0# pfet w=20 l=2
+  ad=240 pd=104 as=320 ps=152
M1001 vdd C out w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 out B vdd w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 vdd A out w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 a_13_n78# D gnd Gnd nfet w=40 l=2
+  ad=240 pd=92 as=200 ps=90
M1005 a_21_n78# C a_13_n78# Gnd nfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1006 a_29_n78# B a_21_n78# Gnd nfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1007 out A a_29_n78# Gnd nfet w=40 l=2
+  ad=280 pd=94 as=0 ps=0
C0 w_0_0# gnd! 1.9fF
