magic
tech scmos
timestamp 1619598226
<< nwell >>
rect 7 77 11 80
rect 38 -91 72 -90
rect 41 -94 72 -91
<< metal1 >>
rect 16 89 63 93
rect -3 80 1 83
rect 16 80 20 89
rect 30 80 34 83
rect 7 77 11 80
rect 59 66 63 89
rect -9 37 4 41
rect -21 30 18 34
rect 25 33 50 34
rect 25 30 57 33
rect 49 29 50 30
rect 72 23 86 27
rect 0 0 74 3
rect -5 -3 74 0
rect 2 -9 26 -3
rect 81 -27 86 23
rect 2 -31 12 -27
rect 30 -33 48 -29
rect 63 -31 86 -27
rect 19 -37 34 -33
rect 71 -38 89 -34
rect 26 -72 32 -70
rect 24 -75 32 -72
rect 28 -91 32 -75
rect 28 -94 40 -91
rect 41 -94 72 -91
<< m2contact >>
rect -14 37 -9 42
rect -26 30 -21 35
rect 89 -38 94 -33
<< metal2 >>
rect -26 35 -21 105
rect -14 42 -9 105
rect 89 -33 94 -11
use 2NAND_WO  2NAND_WO_0
timestamp 1619444932
transform 1 0 1 0 1 50
box -1 -50 32 33
use 2INV  2INV_0
timestamp 1619542334
transform 1 0 50 0 1 -45
box 0 45 24 116
use 2INV  2INV_1
timestamp 1619542334
transform -1 0 26 0 -1 41
box 0 45 24 116
use 2NOR_WO  2NOR_WO_0
timestamp 1619593969
transform -1 0 72 0 -1 -42
box -1 -42 34 52
<< labels >>
rlabel metal2 -12 100 -12 100 5 g1
rlabel metal2 93 -16 93 -16 7 g2
rlabel metal1 36 -93 36 -93 1 gnd
rlabel metal1 42 92 42 92 1 vdd
rlabel metal1 82 25 82 25 1 term1
rlabel metal2 -24 100 -24 100 4 p2
rlabel metal1 38 32 38 32 1 term1_bar
rlabel metal1 24 -35 24 -35 1 out_bar
rlabel metal1 4 -29 4 -29 1 out
<< end >>
