* SPICE3 file created from 3AND.ext - technology: scmos
.option scale=0.09u
.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.global gnd vdd

Vdd	vdd	gnd	'SUPPLY'
vdA     A     0 pulse 1.8 0 0ns 100ps 100ps 5ns  30ns
vdB     B     0 pulse 1.8 0 30ns 100ps 100ps 10ns  30ns

M1000 out_bar out vdd w_51_0# CMOSP w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1001 out_bar out gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=150 ps=90
M1002 a_13_5# B vdd w_0_n1# CMOSP w=40 l=2
+  ad=240 pd=92 as=200 ps=90
M1003 out A a_13_5# w_0_n1# CMOSP w=40 l=2
+  ad=280 pd=94 as=0 ps=0
M1004 out B gnd gnd CMOSN w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1005 gnd A out gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
C0 w_0_n1# gnd 1.9fF




.tran 1n 60n
.control
set hcopypscolor = 1
set color0=white
set color1=black

run
plot v(A) v(B)+2 v(out)+4 v(out_bar)+6
set curplottitle= "Aravind Narayanan-2019102014"
.endc