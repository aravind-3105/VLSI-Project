magic
tech scmos
timestamp 1619522121
<< nwell >>
rect 0 0 41 32
<< ntransistor >>
rect 11 -61 13 -31
rect 19 -61 21 -31
rect 27 -61 29 -31
<< ptransistor >>
rect 11 6 13 26
rect 19 6 21 26
rect 27 6 29 26
<< ndiffusion >>
rect 10 -61 11 -31
rect 13 -61 19 -31
rect 21 -61 27 -31
rect 29 -61 32 -31
<< pdiffusion >>
rect 10 6 11 26
rect 13 6 14 26
rect 18 6 19 26
rect 21 6 22 26
rect 26 6 27 26
rect 29 6 30 26
<< ndcontact >>
rect 6 -61 10 -31
rect 32 -61 36 -31
<< pdcontact >>
rect 6 6 10 26
rect 14 6 18 26
rect 22 6 26 26
rect 30 6 34 26
<< polysilicon >>
rect 11 26 13 29
rect 19 26 21 29
rect 27 26 29 29
rect 11 -24 13 6
rect 19 -17 21 6
rect 27 -10 29 6
rect 11 -31 13 -28
rect 19 -31 21 -21
rect 27 -31 29 -14
rect 11 -64 13 -61
rect 19 -64 21 -61
rect 27 -64 29 -61
<< polycontact >>
rect 25 -14 29 -10
rect 17 -21 21 -17
rect 9 -28 13 -24
<< metal1 >>
rect 0 31 41 34
rect 6 26 10 31
rect 22 26 26 31
rect 14 -3 18 6
rect 30 -3 34 6
rect 14 -7 36 -3
rect 0 -14 25 -10
rect 32 -15 36 -7
rect 0 -21 17 -17
rect 32 -19 41 -15
rect 0 -28 9 -24
rect 32 -31 36 -19
rect 6 -65 10 -61
rect 0 -68 41 -65
<< labels >>
rlabel metal1 7 -12 7 -12 1 A
rlabel metal1 7 -19 7 -19 1 B
rlabel metal1 7 -26 7 -26 1 C
rlabel metal1 39 -17 39 -17 7 out
rlabel metal1 17 33 17 33 5 vdd
rlabel metal1 23 -66 23 -66 1 gnd
<< end >>
