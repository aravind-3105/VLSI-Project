.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.param width_N={10*LAMBDA}
.param width_P={20*LAMBDA}
.global gnd vdd

Vdd	vdd	gnd	'SUPPLY'
vd1a a1  0 pulse 1.8 0 0ns 100ps 100ps 20ns  40ns
vd2a a2  0 pulse 0 0 0ns 100ps 100ps 40ns  80ns
vd3a a3  0 pulse 0 0 0ns 100ps 100ps 80ns  160ns
vd4a a4  0 pulse 0 0 0ns 100ps 100ps 160ns 320ns

vd1b b1  0 pulse 1.8 0 0ns 100ps 100ps 20ns  40ns
vd2b b2  0 pulse 0 0 0ns 100ps 100ps 40ns  80ns
vd3b b3  0 pulse 0 0 0ns 100ps 100ps 80ns  160ns
vd4b b4  0 pulse 0 0 0ns 100ps 100ps 160ns 320ns

M1000 SUM_WO_0/XOR_WO_3/a_59_n30# c4 SUM_WO_0/XOR_WO_3/2INV_1/a_6_87# SUM_WO_0/XOR_WO_3/2INV_1/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1001 SUM_WO_0/XOR_WO_3/a_59_n30# c4 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=3640 ps=2028
M1002 SUM_WO_0/XOR_WO_3/a_51_n59# p4 vdd SUM_WO_0/XOR_WO_3/2INV_0/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=5780 ps=2582
M1003 SUM_WO_0/XOR_WO_3/a_51_n59# p4 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1004 vdd SUM_WO_0/XOR_WO_3/a_51_n59# SUM_WO_0/XOR_WO_3/a_56_27# SUM_WO_0/XOR_WO_3/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=400 ps=180
M1005 SUM_WO_0/XOR_WO_3/a_71_27# SUM_WO_0/XOR_WO_3/a_59_n30# vdd SUM_WO_0/XOR_WO_3/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1006 s4 p4 SUM_WO_0/XOR_WO_3/a_71_27# SUM_WO_0/XOR_WO_3/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1007 SUM_WO_0/XOR_WO_3/a_56_27# c4 s4 SUM_WO_0/XOR_WO_3/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1008 SUM_WO_0/XOR_WO_3/a_63_n51# SUM_WO_0/XOR_WO_3/a_59_n30# gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1009 s4 SUM_WO_0/XOR_WO_3/a_51_n59# SUM_WO_0/XOR_WO_3/a_63_n51# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1010 SUM_WO_0/XOR_WO_3/a_79_n51# p4 s4 Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1011 gnd c4 SUM_WO_0/XOR_WO_3/a_79_n51# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1012 SUM_WO_0/XOR_WO_2/a_59_n30# c3 SUM_WO_0/XOR_WO_2/2INV_1/a_6_87# SUM_WO_0/XOR_WO_2/2INV_1/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1013 SUM_WO_0/XOR_WO_2/a_59_n30# c3 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1014 SUM_WO_0/XOR_WO_2/a_51_n59# p3 vdd SUM_WO_0/XOR_WO_2/2INV_0/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1015 SUM_WO_0/XOR_WO_2/a_51_n59# p3 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1016 vdd SUM_WO_0/XOR_WO_2/a_51_n59# SUM_WO_0/XOR_WO_2/a_56_27# SUM_WO_0/XOR_WO_2/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=400 ps=180
M1017 SUM_WO_0/XOR_WO_2/a_71_27# SUM_WO_0/XOR_WO_2/a_59_n30# vdd SUM_WO_0/XOR_WO_2/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1018 s3 p3 SUM_WO_0/XOR_WO_2/a_71_27# SUM_WO_0/XOR_WO_2/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1019 SUM_WO_0/XOR_WO_2/a_56_27# c3 s3 SUM_WO_0/XOR_WO_2/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1020 SUM_WO_0/XOR_WO_2/a_63_n51# SUM_WO_0/XOR_WO_2/a_59_n30# gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1021 s3 SUM_WO_0/XOR_WO_2/a_51_n59# SUM_WO_0/XOR_WO_2/a_63_n51# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1022 SUM_WO_0/XOR_WO_2/a_79_n51# p3 s3 Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1023 gnd c3 SUM_WO_0/XOR_WO_2/a_79_n51# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1024 SUM_WO_0/XOR_WO_1/a_59_n30# c2 SUM_WO_0/XOR_WO_1/2INV_1/a_6_87# SUM_WO_0/XOR_WO_1/2INV_1/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1025 SUM_WO_0/XOR_WO_1/a_59_n30# c2 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1026 SUM_WO_0/XOR_WO_1/a_51_n59# p2 vdd SUM_WO_0/XOR_WO_1/2INV_0/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1027 SUM_WO_0/XOR_WO_1/a_51_n59# p2 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1028 vdd SUM_WO_0/XOR_WO_1/a_51_n59# SUM_WO_0/XOR_WO_1/a_56_27# SUM_WO_0/XOR_WO_1/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=400 ps=180
M1029 SUM_WO_0/XOR_WO_1/a_71_27# SUM_WO_0/XOR_WO_1/a_59_n30# vdd SUM_WO_0/XOR_WO_1/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1030 s2 p2 SUM_WO_0/XOR_WO_1/a_71_27# SUM_WO_0/XOR_WO_1/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1031 SUM_WO_0/XOR_WO_1/a_56_27# c2 s2 SUM_WO_0/XOR_WO_1/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1032 SUM_WO_0/XOR_WO_1/a_63_n51# SUM_WO_0/XOR_WO_1/a_59_n30# gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1033 s2 SUM_WO_0/XOR_WO_1/a_51_n59# SUM_WO_0/XOR_WO_1/a_63_n51# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1034 SUM_WO_0/XOR_WO_1/a_79_n51# p2 s2 Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1035 gnd c2 SUM_WO_0/XOR_WO_1/a_79_n51# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1036 SUM_WO_0/XOR_WO_0/a_59_n30# g1 SUM_WO_0/XOR_WO_0/2INV_1/a_6_87# SUM_WO_0/XOR_WO_0/2INV_1/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1037 SUM_WO_0/XOR_WO_0/a_59_n30# g1 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1038 SUM_WO_0/XOR_WO_0/a_51_n59# p1 vdd SUM_WO_0/XOR_WO_0/2INV_0/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1039 SUM_WO_0/XOR_WO_0/a_51_n59# p1 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1040 vdd SUM_WO_0/XOR_WO_0/a_51_n59# SUM_WO_0/XOR_WO_0/a_56_27# SUM_WO_0/XOR_WO_0/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=400 ps=180
M1041 SUM_WO_0/XOR_WO_0/a_71_27# SUM_WO_0/XOR_WO_0/a_59_n30# vdd SUM_WO_0/XOR_WO_0/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1042 s1 p1 SUM_WO_0/XOR_WO_0/a_71_27# SUM_WO_0/XOR_WO_0/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1043 SUM_WO_0/XOR_WO_0/a_56_27# g1 s1 SUM_WO_0/XOR_WO_0/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1044 SUM_WO_0/XOR_WO_0/a_63_n51# SUM_WO_0/XOR_WO_0/a_59_n30# gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1045 s1 SUM_WO_0/XOR_WO_0/a_51_n59# SUM_WO_0/XOR_WO_0/a_63_n51# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1046 SUM_WO_0/XOR_WO_0/a_79_n51# p1 s1 Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1047 gnd g1 SUM_WO_0/XOR_WO_0/a_79_n51# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1048 c4 Carry_WO_0/m1_409_n151# Carry_WO_0/2INV_8/a_6_87# Carry_WO_0/2INV_8/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1049 c4 Carry_WO_0/m1_409_n151# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1050 Carry_WO_0/4NOR_WO_0/a_13_6# Carry_WO_0/m1_395_n85# vdd Carry_WO_0/4NOR_WO_0/w_0_0# pfet w=80 l=2
+  ad=480 pd=172 as=0 ps=0
M1051 Carry_WO_0/4NOR_WO_0/a_21_6# Carry_WO_0/m1_402_n83# Carry_WO_0/4NOR_WO_0/a_13_6# Carry_WO_0/4NOR_WO_0/w_0_0# pfet w=80 l=2
+  ad=480 pd=172 as=0 ps=0
M1052 Carry_WO_0/4NOR_WO_0/a_29_6# Carry_WO_0/m1_409_n82# Carry_WO_0/4NOR_WO_0/a_21_6# Carry_WO_0/4NOR_WO_0/w_0_0# pfet w=80 l=2
+  ad=480 pd=172 as=0 ps=0
M1053 Carry_WO_0/m1_409_n151# g4 Carry_WO_0/4NOR_WO_0/a_29_6# Carry_WO_0/4NOR_WO_0/w_0_0# pfet w=80 l=2
+  ad=560 pd=174 as=0 ps=0
M1054 Carry_WO_0/m1_409_n151# Carry_WO_0/m1_395_n85# gnd Gnd nfet w=10 l=2
+  ad=120 pd=64 as=0 ps=0
M1055 gnd Carry_WO_0/m1_402_n83# Carry_WO_0/m1_409_n151# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1056 Carry_WO_0/m1_409_n151# Carry_WO_0/m1_409_n82# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1057 gnd g4 Carry_WO_0/m1_409_n151# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1058 Carry_WO_0/m1_409_n82# Carry_WO_0/m1_683_20# Carry_WO_0/2INV_7/a_6_87# Carry_WO_0/2INV_7/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1059 Carry_WO_0/m1_409_n82# Carry_WO_0/m1_683_20# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1060 Carry_WO_0/m1_683_20# p4 vdd Carry_WO_0/4NAND_WO_0/w_0_0# pfet w=20 l=2
+  ad=240 pd=104 as=0 ps=0
M1061 vdd p3 Carry_WO_0/m1_683_20# Carry_WO_0/4NAND_WO_0/w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1062 Carry_WO_0/m1_683_20# p2 vdd Carry_WO_0/4NAND_WO_0/w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1063 vdd g1 Carry_WO_0/m1_683_20# Carry_WO_0/4NAND_WO_0/w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1064 Carry_WO_0/4NAND_WO_0/a_13_n78# p4 gnd Gnd nfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1065 Carry_WO_0/4NAND_WO_0/a_21_n78# p3 Carry_WO_0/4NAND_WO_0/a_13_n78# Gnd nfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1066 Carry_WO_0/4NAND_WO_0/a_29_n78# p2 Carry_WO_0/4NAND_WO_0/a_21_n78# Gnd nfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1067 Carry_WO_0/m1_683_20# g1 Carry_WO_0/4NAND_WO_0/a_29_n78# Gnd nfet w=40 l=2
+  ad=280 pd=94 as=0 ps=0
M1068 Carry_WO_0/3NOR_WO_0/a_14_3# Carry_WO_0/m1_174_23# vdd Carry_WO_0/3NOR_WO_0/w_1_n3# pfet w=60 l=2
+  ad=360 pd=132 as=0 ps=0
M1069 Carry_WO_0/3NOR_WO_0/a_22_3# g3 Carry_WO_0/3NOR_WO_0/a_14_3# Carry_WO_0/3NOR_WO_0/w_1_n3# pfet w=60 l=2
+  ad=360 pd=132 as=0 ps=0
M1070 Carry_WO_0/m1_194_n80# Carry_WO_0/m1_226_n94# Carry_WO_0/3NOR_WO_0/a_22_3# Carry_WO_0/3NOR_WO_0/w_1_n3# pfet w=60 l=2
+  ad=420 pd=134 as=0 ps=0
M1071 Carry_WO_0/m1_194_n80# Carry_WO_0/m1_174_23# gnd Gnd nfet w=10 l=2
+  ad=130 pd=66 as=0 ps=0
M1072 gnd g3 Carry_WO_0/m1_194_n80# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1073 Carry_WO_0/m1_194_n80# Carry_WO_0/m1_226_n94# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1074 c3 Carry_WO_0/m1_194_n80# Carry_WO_0/2INV_3/a_6_87# Carry_WO_0/2INV_3/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1075 c3 Carry_WO_0/m1_194_n80# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1076 Carry_WO_0/m1_402_n83# Carry_WO_0/m1_526_53# Carry_WO_0/2INV_6/a_6_87# Carry_WO_0/2INV_6/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1077 Carry_WO_0/m1_402_n83# Carry_WO_0/m1_526_53# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1078 Carry_WO_0/m1_526_53# p4 vdd Carry_WO_0/3NAND_WO_1/w_0_0# pfet w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M1079 vdd p3 Carry_WO_0/m1_526_53# Carry_WO_0/3NAND_WO_1/w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1080 Carry_WO_0/m1_526_53# g2 vdd Carry_WO_0/3NAND_WO_1/w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1081 Carry_WO_0/3NAND_WO_1/a_13_n61# p4 gnd Gnd nfet w=30 l=2
+  ad=180 pd=72 as=0 ps=0
M1082 Carry_WO_0/3NAND_WO_1/a_21_n61# p3 Carry_WO_0/3NAND_WO_1/a_13_n61# Gnd nfet w=30 l=2
+  ad=180 pd=72 as=0 ps=0
M1083 Carry_WO_0/m1_526_53# g2 Carry_WO_0/3NAND_WO_1/a_21_n61# Gnd nfet w=30 l=2
+  ad=210 pd=74 as=0 ps=0
M1084 Carry_WO_0/m1_395_n85# Carry_WO_0/m1_398_36# Carry_WO_0/2INV_5/a_6_87# Carry_WO_0/2INV_5/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1085 Carry_WO_0/m1_395_n85# Carry_WO_0/m1_398_36# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1086 Carry_WO_0/m1_398_36# p4 vdd Carry_WO_0/2NAND_WO_2/w_0_0# pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1087 vdd g3 Carry_WO_0/m1_398_36# Carry_WO_0/2NAND_WO_2/w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1088 Carry_WO_0/2NAND_WO_2/a_13_n43# p4 gnd Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1089 Carry_WO_0/m1_398_36# g3 Carry_WO_0/2NAND_WO_2/a_13_n43# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1090 Carry_WO_0/m1_226_n94# Carry_WO_0/m1_252_46# Carry_WO_0/2INV_4/a_6_87# Carry_WO_0/2INV_4/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1091 Carry_WO_0/m1_226_n94# Carry_WO_0/m1_252_46# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1092 Carry_WO_0/m1_252_46# g1 vdd Carry_WO_0/3NAND_WO_0/w_0_0# pfet w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M1093 vdd p2 Carry_WO_0/m1_252_46# Carry_WO_0/3NAND_WO_0/w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1094 Carry_WO_0/m1_252_46# p3 vdd Carry_WO_0/3NAND_WO_0/w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1095 Carry_WO_0/3NAND_WO_0/a_13_n61# g1 gnd Gnd nfet w=30 l=2
+  ad=180 pd=72 as=0 ps=0
M1096 Carry_WO_0/3NAND_WO_0/a_21_n61# p2 Carry_WO_0/3NAND_WO_0/a_13_n61# Gnd nfet w=30 l=2
+  ad=180 pd=72 as=0 ps=0
M1097 Carry_WO_0/m1_252_46# p3 Carry_WO_0/3NAND_WO_0/a_21_n61# Gnd nfet w=30 l=2
+  ad=210 pd=74 as=0 ps=0
M1098 Carry_WO_0/m1_174_23# Carry_WO_0/m1_145_29# Carry_WO_0/2INV_2/a_6_87# Carry_WO_0/2INV_2/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1099 Carry_WO_0/m1_174_23# Carry_WO_0/m1_145_29# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1100 Carry_WO_0/m1_145_29# p3 vdd Carry_WO_0/2NAND_WO_1/w_0_0# pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1101 vdd g2 Carry_WO_0/m1_145_29# Carry_WO_0/2NAND_WO_1/w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1102 Carry_WO_0/2NAND_WO_1/a_13_n43# p3 gnd Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1103 Carry_WO_0/m1_145_29# g2 Carry_WO_0/2NAND_WO_1/a_13_n43# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1104 Carry_WO_0/2NOR_WO_0/a_13_5# Carry_WO_0/m1_63_n31# vdd Carry_WO_0/w_38_n91# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1105 Carry_WO_0/m1_19_n37# g2 Carry_WO_0/2NOR_WO_0/a_13_5# Carry_WO_0/w_38_n91# pfet w=40 l=2
+  ad=280 pd=94 as=0 ps=0
M1106 Carry_WO_0/m1_19_n37# Carry_WO_0/m1_63_n31# gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1107 gnd g2 Carry_WO_0/m1_19_n37# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1108 c2 Carry_WO_0/m1_19_n37# Carry_WO_0/2INV_1/a_6_87# Carry_WO_0/2INV_1/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1109 c2 Carry_WO_0/m1_19_n37# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1110 Carry_WO_0/m1_63_n31# Carry_WO_0/m1_25_30# Carry_WO_0/2INV_0/a_6_87# Carry_WO_0/2INV_0/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1111 Carry_WO_0/m1_63_n31# Carry_WO_0/m1_25_30# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1112 Carry_WO_0/m1_25_30# g1 vdd Carry_WO_0/w_7_77# pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1113 vdd p2 Carry_WO_0/m1_25_30# Carry_WO_0/w_7_77# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1114 Carry_WO_0/2NAND_WO_0/a_13_n43# g1 gnd Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1115 Carry_WO_0/m1_25_30# p2 Carry_WO_0/2NAND_WO_0/a_13_n43# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1116 PropGen_WO_0/XOR_WO_3/a_59_n30# b3 PropGen_WO_0/XOR_WO_3/2INV_1/a_6_87# PropGen_WO_0/XOR_WO_3/2INV_1/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1117 PropGen_WO_0/XOR_WO_3/a_59_n30# b3 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1118 PropGen_WO_0/XOR_WO_3/a_51_n59# a3 vdd PropGen_WO_0/XOR_WO_3/2INV_0/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1119 PropGen_WO_0/XOR_WO_3/a_51_n59# a3 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1120 vdd PropGen_WO_0/XOR_WO_3/a_51_n59# PropGen_WO_0/XOR_WO_3/a_56_27# PropGen_WO_0/XOR_WO_3/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=400 ps=180
M1121 PropGen_WO_0/XOR_WO_3/a_71_27# PropGen_WO_0/XOR_WO_3/a_59_n30# vdd PropGen_WO_0/XOR_WO_3/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1122 p4 a3 PropGen_WO_0/XOR_WO_3/a_71_27# PropGen_WO_0/XOR_WO_3/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1123 PropGen_WO_0/XOR_WO_3/a_56_27# b3 p4 PropGen_WO_0/XOR_WO_3/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1124 PropGen_WO_0/XOR_WO_3/a_63_n51# PropGen_WO_0/XOR_WO_3/a_59_n30# gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1125 p4 PropGen_WO_0/XOR_WO_3/a_51_n59# PropGen_WO_0/XOR_WO_3/a_63_n51# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1126 PropGen_WO_0/XOR_WO_3/a_79_n51# a3 p4 Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1127 gnd b3 PropGen_WO_0/XOR_WO_3/a_79_n51# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1128 PropGen_WO_0/XOR_WO_2/a_59_n30# b2 PropGen_WO_0/XOR_WO_2/2INV_1/a_6_87# PropGen_WO_0/XOR_WO_2/2INV_1/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1129 PropGen_WO_0/XOR_WO_2/a_59_n30# b2 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1130 PropGen_WO_0/XOR_WO_2/a_51_n59# a2 vdd PropGen_WO_0/XOR_WO_2/2INV_0/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1131 PropGen_WO_0/XOR_WO_2/a_51_n59# a2 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1132 vdd PropGen_WO_0/XOR_WO_2/a_51_n59# PropGen_WO_0/XOR_WO_2/a_56_27# PropGen_WO_0/XOR_WO_2/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=400 ps=180
M1133 PropGen_WO_0/XOR_WO_2/a_71_27# PropGen_WO_0/XOR_WO_2/a_59_n30# vdd PropGen_WO_0/XOR_WO_2/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1134 p3 a2 PropGen_WO_0/XOR_WO_2/a_71_27# PropGen_WO_0/XOR_WO_2/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1135 PropGen_WO_0/XOR_WO_2/a_56_27# b2 p3 PropGen_WO_0/XOR_WO_2/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1136 PropGen_WO_0/XOR_WO_2/a_63_n51# PropGen_WO_0/XOR_WO_2/a_59_n30# gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1137 p3 PropGen_WO_0/XOR_WO_2/a_51_n59# PropGen_WO_0/XOR_WO_2/a_63_n51# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1138 PropGen_WO_0/XOR_WO_2/a_79_n51# a2 p3 Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1139 gnd b2 PropGen_WO_0/XOR_WO_2/a_79_n51# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1140 PropGen_WO_0/XOR_WO_1/a_59_n30# b1 PropGen_WO_0/XOR_WO_1/2INV_1/a_6_87# PropGen_WO_0/XOR_WO_1/2INV_1/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1141 PropGen_WO_0/XOR_WO_1/a_59_n30# b1 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1142 PropGen_WO_0/XOR_WO_1/a_51_n59# a1 vdd PropGen_WO_0/XOR_WO_1/2INV_0/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1143 PropGen_WO_0/XOR_WO_1/a_51_n59# a1 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1144 vdd PropGen_WO_0/XOR_WO_1/a_51_n59# PropGen_WO_0/XOR_WO_1/a_56_27# PropGen_WO_0/XOR_WO_1/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=400 ps=180
M1145 PropGen_WO_0/XOR_WO_1/a_71_27# PropGen_WO_0/XOR_WO_1/a_59_n30# vdd PropGen_WO_0/XOR_WO_1/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1146 p2 a1 PropGen_WO_0/XOR_WO_1/a_71_27# PropGen_WO_0/XOR_WO_1/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1147 PropGen_WO_0/XOR_WO_1/a_56_27# b1 p2 PropGen_WO_0/XOR_WO_1/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1148 PropGen_WO_0/XOR_WO_1/a_63_n51# PropGen_WO_0/XOR_WO_1/a_59_n30# gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1149 p2 PropGen_WO_0/XOR_WO_1/a_51_n59# PropGen_WO_0/XOR_WO_1/a_63_n51# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1150 PropGen_WO_0/XOR_WO_1/a_79_n51# a1 p2 Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1151 gnd b1 PropGen_WO_0/XOR_WO_1/a_79_n51# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1152 PropGen_WO_0/XOR_WO_0/a_59_n30# b0 PropGen_WO_0/XOR_WO_0/2INV_1/a_6_87# PropGen_WO_0/XOR_WO_0/2INV_1/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1153 PropGen_WO_0/XOR_WO_0/a_59_n30# b0 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1154 PropGen_WO_0/XOR_WO_0/a_51_n59# a0 vdd PropGen_WO_0/XOR_WO_0/2INV_0/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1155 PropGen_WO_0/XOR_WO_0/a_51_n59# a0 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1156 vdd PropGen_WO_0/XOR_WO_0/a_51_n59# PropGen_WO_0/XOR_WO_0/a_56_27# PropGen_WO_0/XOR_WO_0/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=400 ps=180
M1157 PropGen_WO_0/XOR_WO_0/a_71_27# PropGen_WO_0/XOR_WO_0/a_59_n30# vdd PropGen_WO_0/XOR_WO_0/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1158 p1 a0 PropGen_WO_0/XOR_WO_0/a_71_27# PropGen_WO_0/XOR_WO_0/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1159 PropGen_WO_0/XOR_WO_0/a_56_27# b0 p1 PropGen_WO_0/XOR_WO_0/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1160 PropGen_WO_0/XOR_WO_0/a_63_n51# PropGen_WO_0/XOR_WO_0/a_59_n30# gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1161 p1 PropGen_WO_0/XOR_WO_0/a_51_n59# PropGen_WO_0/XOR_WO_0/a_63_n51# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1162 PropGen_WO_0/XOR_WO_0/a_79_n51# a0 p1 Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1163 gnd b0 PropGen_WO_0/XOR_WO_0/a_79_n51# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1164 g2 a1 vdd PropGen_WO_0/2AND_WO_1/w_0_0# pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1165 vdd b1 g2 PropGen_WO_0/2AND_WO_1/w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1166 PropGen_WO_0/2AND_WO_1/a_13_n43# a1 gnd Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1167 g2 b1 PropGen_WO_0/2AND_WO_1/a_13_n43# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1168 g4 a3 vdd PropGen_WO_0/2AND_WO_3/w_0_0# pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1169 vdd b3 g4 PropGen_WO_0/2AND_WO_3/w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1170 PropGen_WO_0/2AND_WO_3/a_13_n43# a3 gnd Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1171 g4 b3 PropGen_WO_0/2AND_WO_3/a_13_n43# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1172 g1 a0 vdd PropGen_WO_0/2AND_WO_0/w_0_0# pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1173 vdd b0 g1 PropGen_WO_0/2AND_WO_0/w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1174 PropGen_WO_0/2AND_WO_0/a_13_n43# a0 gnd Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1175 g1 b0 PropGen_WO_0/2AND_WO_0/a_13_n43# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1176 g3 a2 vdd PropGen_WO_0/2AND_WO_2/w_0_0# pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1177 vdd b2 g3 PropGen_WO_0/2AND_WO_2/w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1178 PropGen_WO_0/2AND_WO_2/a_13_n43# a2 gnd Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1179 g3 b2 PropGen_WO_0/2AND_WO_2/a_13_n43# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
C0 p2 g1 8.3fF
C1 Carry_WO_0/m1_409_n82# Carry_WO_0/m1_402_n83# 2.3fF
C2 g1 vdd 1.9fF
C3 g4 g3 2.0fF
C4 g1 p1 2.8fF
C5 a1 b1 4.8fF
C6 c4 p4 2.0fF
C7 g2 Carry_WO_0/m1_63_n31# 1.2fF
C8 SUM_WO_0/XOR_WO_3/a_56_27# s4 1.1fF
C9 c2 p2 2.0fF
C10 p4 p3 4.3fF
C11 p4 g3 2.9fF
C12 Carry_WO_0/m1_402_n83# Carry_WO_0/m1_395_n85# 1.5fF
C13 a3 b2 5.2fF
C14 a2 b1 2.4fF
C15 g2 p3 6.4fF
C16 g3 p3 2.1fF
C17 c3 p3 2.1fF
C18 a0 b0 3.5fF
C19 SUM_WO_0/XOR_WO_2/a_56_27# s3 1.1fF
C20 p4 PropGen_WO_0/XOR_WO_3/a_56_27# 1.1fF
C21 a2 b2 7.6fF
C22 SUM_WO_0/XOR_WO_0/a_56_27# s1 1.1fF
C23 PropGen_WO_0/XOR_WO_0/a_56_27# p1 1.1fF
C24 SUM_WO_0/XOR_WO_1/a_56_27# s2 1.1fF
C25 g4 Carry_WO_0/m1_409_n82# 2.9fF
C26 p2 p3 4.7fF
C27 p2 g2 2.5fF
C28 vdd p3 1.1fF
C29 g4 p4 2.0fF
C30 p2 PropGen_WO_0/XOR_WO_1/a_56_27# 1.1fF
C31 p3 PropGen_WO_0/XOR_WO_2/a_56_27# 1.1fF
C32 g3 Carry_WO_0/m1_226_n94# 1.1fF
C33 a3 b3 12.8fF
C34 b2 gnd! 5.3fF
C35 PropGen_WO_0/2AND_WO_2/w_0_0# gnd! 1.0fF
C36 b0 gnd! 3.8fF
C37 PropGen_WO_0/2AND_WO_0/w_0_0# gnd! 1.0fF
C38 PropGen_WO_0/2AND_WO_3/w_0_0# gnd! 1.0fF
C39 PropGen_WO_0/2AND_WO_1/w_0_0# gnd! 1.0fF
C40 p1 gnd! 19.6fF
C41 PropGen_WO_0/XOR_WO_0/w_50_21# gnd! 2.7fF
C42 PropGen_WO_0/XOR_WO_0/a_51_n59# gnd! 1.6fF
C43 a0 gnd! 3.8fF
C44 PropGen_WO_0/XOR_WO_1/w_50_21# gnd! 2.7fF
C45 PropGen_WO_0/XOR_WO_1/a_51_n59# gnd! 1.6fF
C46 a1 gnd! 4.3fF
C47 b1 gnd! 5.1fF
C48 p3 gnd! 25.8fF
C49 PropGen_WO_0/XOR_WO_2/w_50_21# gnd! 2.7fF
C50 PropGen_WO_0/XOR_WO_2/a_51_n59# gnd! 1.6fF
C51 a2 gnd! 4.9fF
C52 p4 gnd! 24.5fF
C53 PropGen_WO_0/XOR_WO_3/w_50_21# gnd! 2.7fF
C54 PropGen_WO_0/XOR_WO_3/a_51_n59# gnd! 1.6fF
C55 a3 gnd! 6.9fF
C56 b3 gnd! 6.8fF
C57 Carry_WO_0/w_7_77# gnd! 1.0fF
C58 Carry_WO_0/w_38_n91# gnd! 1.8fF
C59 Carry_WO_0/2NAND_WO_1/w_0_0# gnd! 1.0fF
C60 Carry_WO_0/m1_174_23# gnd! 1.2fF
C61 Carry_WO_0/3NAND_WO_0/w_0_0# gnd! 1.3fF
C62 g3 gnd! 15.3fF
C63 Carry_WO_0/2NAND_WO_2/w_0_0# gnd! 1.0fF
C64 Carry_WO_0/m1_395_n85# gnd! 1.5fF
C65 g2 gnd! 15.1fF
C66 Carry_WO_0/3NAND_WO_1/w_0_0# gnd! 1.3fF
C67 vdd gnd! 55.6fF
C68 Carry_WO_0/m1_402_n83# gnd! 1.9fF
C69 Carry_WO_0/3NOR_WO_0/w_1_n3# gnd! 3.1fF
C70 g1 gnd! 19.7fF
C71 p2 gnd! 24.8fF
C72 Carry_WO_0/4NAND_WO_0/w_0_0# gnd! 1.7fF
C73 gnd gnd! 50.4fF
C74 Carry_WO_0/m1_409_n82# gnd! 4.6fF
C75 g4 gnd! 15.3fF
C76 Carry_WO_0/4NOR_WO_0/w_0_0# gnd! 4.6fF
C77 s1 gnd! 1.5fF
C78 SUM_WO_0/XOR_WO_0/w_50_21# gnd! 2.7fF
C79 SUM_WO_0/XOR_WO_0/a_51_n59# gnd! 1.6fF
C80 s2 gnd! 1.5fF
C81 SUM_WO_0/XOR_WO_1/w_50_21# gnd! 2.7fF
C82 SUM_WO_0/XOR_WO_1/a_51_n59# gnd! 1.6fF
C83 c2 gnd! 7.3fF
C84 s3 gnd! 1.5fF
C85 SUM_WO_0/XOR_WO_2/w_50_21# gnd! 2.7fF
C86 SUM_WO_0/XOR_WO_2/a_51_n59# gnd! 1.6fF
C87 c3 gnd! 6.5fF
C88 s4 gnd! 1.6fF
C89 SUM_WO_0/XOR_WO_3/w_50_21# gnd! 2.7fF
C90 SUM_WO_0/XOR_WO_3/a_51_n59# gnd! 1.6fF
C91 c4 gnd! 5.9fF



.ic v(a1) = 0
.ic v(b1) = 0
.ic v(a2) = 0
.ic v(b2) = 0
.ic v(a3) = 0
.ic v(b3) = 0
.ic v(a4) = 0
.ic v(b4) = 0
.tran 0.01n 40n
.control
set hcopypscolor = 1
set color0=white
set color1=black

run
plot v(a1)/1.8 ((v(b1)/1.8)+4)
plot v(a2)/1.8 ((v(b2)/1.8)+4)
plot v(a3)/1.8 ((v(b3)/1.8)+4)
plot v(a4)/1.8 ((v(b4)/1.8)+4)
plot (v(a1)+(2*v(a2))+(4*v(a3))+(8*v(a4)))/1.8
plot (v(b1)+(2*v(b2))+(4*v(b3))+(8*v(b4)))/1.8
* plot (v(Sum1)+(2*v(Sum2))+(4*v(Sum3))+(8*v(Sum4)))/1.8
* plot v(Cout4)/1.8
set curplottitle= "Aravind Narayanan-2019102014"
.endc