magic
tech scmos
timestamp 1619686085
<< metal1 >>
rect -201 820 -177 824
rect -171 820 -14 824
rect -362 760 -341 764
rect -188 758 -120 762
rect -419 605 -414 751
rect -419 542 -414 600
rect -432 534 -414 542
rect -419 453 -414 534
rect -419 299 -414 448
rect -419 147 -414 294
rect -419 -8 -414 141
rect -419 -244 -414 -14
rect -377 703 -334 707
rect -377 559 -371 703
rect -124 692 -120 758
rect -18 744 -14 820
rect -18 740 19 744
rect 21 701 26 731
rect 87 707 92 734
rect 113 701 118 731
rect 179 713 184 743
rect 1842 738 1849 740
rect 1842 734 2023 738
rect -185 671 -177 675
rect -346 611 -336 615
rect -114 613 -109 678
rect -185 609 -109 613
rect 1473 671 1758 678
rect -354 606 -349 608
rect 325 604 526 609
rect -377 554 -335 559
rect 21 556 26 586
rect 87 562 92 589
rect 113 556 118 586
rect 179 563 184 593
rect -377 409 -371 554
rect -189 521 -177 525
rect -106 463 -101 542
rect -193 459 -101 463
rect -351 454 -348 458
rect -95 453 -89 533
rect -163 449 -89 453
rect -377 404 -335 409
rect -377 258 -371 404
rect -163 312 -157 449
rect 21 411 26 441
rect 87 417 92 444
rect 113 411 118 441
rect 179 420 184 450
rect -188 308 -157 312
rect -352 300 -348 307
rect -124 272 -118 397
rect -167 267 -118 272
rect -377 253 -335 258
rect -377 107 -371 253
rect -192 219 -177 223
rect -167 161 -164 267
rect -108 262 -103 384
rect 205 342 237 347
rect 195 305 212 309
rect 240 299 289 303
rect 21 265 26 295
rect 113 265 118 295
rect -189 157 -164 161
rect -159 258 -103 262
rect 205 259 237 264
rect -353 148 -349 156
rect -377 102 -336 107
rect -377 -44 -371 102
rect -190 68 -177 72
rect -159 35 -153 258
rect -159 10 -154 35
rect -188 6 -154 10
rect -353 -8 -349 5
rect -156 -38 -152 -21
rect -123 -26 -119 247
rect -110 -17 -106 231
rect 201 222 209 226
rect 325 220 329 604
rect 242 219 329 220
rect 219 216 329 219
rect 319 212 329 216
rect 205 155 237 160
rect 359 157 363 561
rect 294 153 363 157
rect 199 103 202 122
rect 240 112 319 116
rect 315 111 319 112
rect 409 111 413 561
rect 315 106 413 111
rect 167 81 237 86
rect 447 54 452 563
rect 603 152 609 230
rect 773 189 778 215
rect 1015 210 1019 231
rect 1473 210 1478 671
rect 1842 666 1849 734
rect 2118 733 2171 737
rect 1945 673 1991 677
rect 1567 657 1849 666
rect 1567 569 1574 657
rect 1735 656 1849 657
rect 1920 666 2009 670
rect 1760 647 1864 652
rect 1760 643 1764 647
rect 1567 564 1591 569
rect 1920 493 1923 666
rect 1968 615 2003 621
rect 2166 564 2171 733
rect 2146 560 2171 564
rect 1944 500 1988 504
rect 1956 493 2009 497
rect 1920 488 1959 493
rect 1761 447 1883 451
rect 1560 406 1565 421
rect 1015 205 1478 210
rect 1522 402 1565 406
rect 1522 189 1527 402
rect 773 184 1527 189
rect 1539 152 1545 354
rect 1920 336 1923 488
rect 1981 443 2001 448
rect 2166 403 2171 560
rect 2146 399 2171 403
rect 1984 339 1988 343
rect 1920 332 1995 336
rect 1760 298 1878 304
rect 1922 183 1928 332
rect 1963 282 1997 287
rect 2166 250 2171 399
rect 2149 246 2171 250
rect 1984 186 1986 190
rect 1922 179 1990 183
rect 603 147 1545 152
rect 243 50 452 54
rect 1395 51 1400 112
rect 195 44 208 48
rect 243 38 246 50
rect 1553 51 1558 147
rect 1760 141 1887 146
rect 307 20 523 23
rect 224 18 523 20
rect 224 15 311 18
rect 1759 -14 1764 71
rect 1922 49 1928 179
rect 1974 130 2002 134
rect 1969 129 2002 130
rect 2166 78 2171 246
rect 2147 74 2171 78
rect -110 -21 58 -17
rect 1921 11 1928 49
rect 1921 7 2007 11
rect -123 -29 -90 -26
rect -94 -37 -90 -29
rect 54 -37 58 -21
rect 586 -39 592 -38
rect 1921 -39 1928 7
rect -377 -49 -341 -44
rect -188 -220 -183 -44
rect 586 -51 1928 -39
rect 1956 -43 2005 -38
rect 111 -143 524 -139
rect -96 -209 -92 -194
rect -89 -198 -85 -197
rect -40 -220 -35 -176
rect 59 -202 63 -195
rect 59 -206 67 -202
rect 108 -220 113 -186
rect -188 -226 113 -220
rect 586 -244 592 -51
rect -419 -254 -66 -244
rect -57 -254 67 -244
rect 74 -253 592 -244
rect 74 -254 86 -253
rect 586 -254 592 -253
<< m2contact >>
rect -177 819 -171 824
rect -368 760 -362 765
rect -419 751 -414 756
rect -353 752 -348 757
rect -419 600 -414 605
rect -419 448 -414 453
rect -419 294 -414 299
rect -419 141 -414 147
rect -419 -14 -414 -8
rect -124 687 -119 692
rect -114 678 -109 683
rect -177 670 -171 675
rect -351 611 -346 616
rect 1758 671 1764 678
rect -354 601 -349 606
rect 526 604 531 609
rect -106 542 -101 547
rect -177 520 -171 525
rect -351 461 -346 466
rect -95 533 -89 538
rect -353 449 -348 454
rect -351 310 -345 315
rect -124 397 -118 402
rect -352 295 -347 300
rect -108 384 -103 389
rect -177 218 -171 223
rect -352 159 -347 164
rect 289 298 294 303
rect -354 142 -348 148
rect -177 67 -171 73
rect -124 247 -119 252
rect -353 8 -348 13
rect -353 -13 -348 -8
rect -157 -21 -152 -16
rect -110 231 -105 236
rect 359 561 364 566
rect 409 561 414 566
rect 447 563 452 568
rect 289 153 294 158
rect 1940 673 1945 678
rect 2150 671 2155 676
rect 1960 615 1968 621
rect 1939 499 1944 505
rect 2149 498 2154 503
rect 1883 447 1889 452
rect 1560 421 1565 426
rect 1539 354 1545 359
rect 1976 443 1981 449
rect 1978 339 1984 344
rect 2150 337 2155 342
rect 1878 298 1883 304
rect 1956 282 1963 287
rect 1978 186 1984 191
rect 1553 147 1558 152
rect 1395 112 1400 117
rect 1395 46 1400 51
rect 1587 137 1592 142
rect 1887 141 1893 146
rect 1553 46 1558 51
rect 523 18 528 23
rect 1968 130 1974 135
rect 1759 -19 1764 -14
rect 1983 14 1988 19
rect 2148 12 2153 17
rect -8 -38 -3 -33
rect 1949 -43 1956 -37
rect 524 -143 529 -137
rect -89 -203 -84 -198
rect -97 -214 -92 -209
rect 67 -206 72 -201
rect -66 -238 -61 -233
rect -66 -254 -57 -244
rect 67 -254 74 -244
<< metal2 >>
rect -423 760 -368 765
rect -414 752 -353 756
rect -177 675 -171 819
rect 301 811 530 814
rect 105 809 530 811
rect 105 807 307 809
rect 185 806 307 807
rect -119 687 -85 692
rect -124 678 -114 683
rect -109 678 -85 683
rect -423 611 -351 615
rect -423 610 -369 611
rect -414 601 -354 605
rect -414 600 -381 601
rect -177 525 -171 670
rect 307 667 474 670
rect 106 665 474 667
rect 106 663 310 665
rect 194 662 310 663
rect 470 638 474 665
rect 526 668 530 809
rect 1764 673 1940 677
rect 2155 671 2181 675
rect 526 663 625 668
rect 1362 663 1554 668
rect 516 653 529 658
rect 493 643 528 648
rect 470 633 723 638
rect 1366 633 1524 638
rect 364 623 590 628
rect 322 613 538 618
rect 1346 613 1500 618
rect -124 542 -106 547
rect -101 542 -85 547
rect -124 533 -95 538
rect -89 533 -85 538
rect 322 527 326 613
rect 1370 604 1395 609
rect 359 566 364 573
rect 409 566 414 573
rect 504 568 509 572
rect 452 564 509 568
rect 189 523 326 527
rect 106 522 326 523
rect 486 535 609 540
rect 106 520 311 522
rect -428 461 -351 465
rect -414 449 -353 453
rect -422 310 -351 314
rect -414 295 -352 299
rect -177 223 -171 520
rect 189 519 311 520
rect -118 397 -95 402
rect -89 397 -85 402
rect -124 384 -108 389
rect -103 384 -96 389
rect -88 384 -63 389
rect 189 372 425 377
rect 189 369 319 372
rect -105 247 -85 252
rect -105 231 -85 236
rect -424 159 -352 163
rect -414 142 -354 147
rect -177 73 -171 218
rect 289 158 294 298
rect 420 129 425 372
rect 486 142 490 535
rect -424 8 -353 12
rect -414 -13 -353 -8
rect -177 -16 -171 67
rect -177 -21 -157 -16
rect -152 -21 -3 -16
rect -8 -33 -3 -21
rect 167 -32 172 4
rect 167 -33 173 -32
rect 486 -33 490 137
rect 524 23 528 467
rect 1496 219 1500 613
rect 1520 368 1524 633
rect 1548 515 1554 663
rect 1859 647 1966 652
rect 1686 634 1943 639
rect 1548 510 1615 515
rect 1939 505 1943 634
rect 1960 621 1966 647
rect 1560 500 1625 505
rect 1560 426 1565 500
rect 2154 498 2190 502
rect 1686 485 1835 490
rect 1520 363 1643 368
rect 1545 354 1579 359
rect 1830 344 1835 485
rect 1889 449 1980 451
rect 1889 447 1976 449
rect 1686 338 1792 343
rect 1830 339 1978 344
rect 1787 231 1792 338
rect 2155 337 2194 341
rect 1883 298 1961 304
rect 1956 287 1961 298
rect 1787 226 1872 231
rect 1496 214 1643 219
rect 1553 205 1577 210
rect 1553 152 1558 205
rect 1686 186 1821 191
rect 1867 190 1872 226
rect 1867 186 1978 190
rect 1984 186 1989 190
rect 563 137 1587 142
rect 538 60 543 124
rect 1395 117 1400 122
rect 538 55 1638 60
rect 1400 46 1553 51
rect 167 -39 490 -33
rect 524 -14 528 18
rect 1575 -14 1582 51
rect 1664 46 1735 51
rect 1816 18 1821 186
rect 2154 184 2185 188
rect 1893 141 1973 146
rect 1968 135 1973 141
rect 1968 129 1973 130
rect 1816 14 1983 18
rect 1988 14 1989 18
rect 2153 12 2188 16
rect 582 -19 1759 -14
rect 1764 -19 1954 -14
rect -426 -71 -256 -66
rect -426 -87 -283 -81
rect -289 -220 -283 -87
rect -262 -209 -256 -71
rect -84 -203 -66 -199
rect -262 -214 -97 -209
rect 52 -220 56 -193
rect -289 -226 56 -220
rect -66 -244 -61 -238
rect 67 -244 71 -206
rect 325 -269 336 -39
rect 524 -137 529 -19
rect 1949 -37 1954 -19
rect 524 -270 529 -143
<< m3contact >>
rect 511 653 516 658
rect 488 643 493 648
rect 359 623 364 628
rect 1395 604 1400 609
rect 359 573 364 578
rect 409 573 414 578
rect 504 572 509 577
rect 420 124 425 129
rect 486 137 491 142
rect 558 137 563 142
rect 538 124 543 129
rect 1395 122 1400 127
rect 524 -19 529 -14
rect 577 -19 582 -14
rect -66 -203 -61 -198
<< metal3 >>
rect 504 653 511 658
rect 409 643 488 648
rect 359 578 364 623
rect 409 578 414 643
rect 504 577 509 653
rect 491 137 558 142
rect 425 124 538 129
rect 1395 127 1400 604
rect 529 -19 577 -14
rect -66 -238 -61 -203
use FlipFlop_WO  FlipFlop_WO_5
timestamp 1619646873
transform 1 0 -349 0 1 767
box -1 -64 165 57
use FlipFlop_WO  FlipFlop_WO_6
timestamp 1619646873
transform 1 0 -349 0 1 618
box -1 -64 165 57
use FlipFlop_WO  FlipFlop_WO_7
timestamp 1619646873
transform 1 0 -350 0 1 468
box -1 -64 165 57
use FlipFlop_WO  FlipFlop_WO_8
timestamp 1619646873
transform 1 0 -351 0 1 317
box -1 -64 165 57
use FlipFlop_WO  FlipFlop_WO_9
timestamp 1619646873
transform 1 0 -352 0 1 166
box -1 -64 165 57
use FlipFlop_WO  FlipFlop_WO_10
timestamp 1619646873
transform 1 0 -352 0 1 15
box -1 -64 165 57
use PropagateGenerate_WO  PropagateGenerate_WO_0
timestamp 1619651442
transform 0 -1 184 1 0 251
box -254 -59 560 308
use Carry_WO  Carry_WO_0
timestamp 1619609411
transform 1 0 612 0 1 455
box -86 -250 759 213
use SUM_WO  SUM_WO_0
timestamp 1619592134
transform 0 -1 1764 1 0 65
box -19 -16 579 189
use FlipFlop_WO  FlipFlop_WO_0
timestamp 1619646873
transform 1 0 1987 0 1 680
box -1 -64 165 57
use FlipFlop_WO  FlipFlop_WO_1
timestamp 1619646873
transform 1 0 1986 0 1 507
box -1 -64 165 57
use FlipFlop_WO  FlipFlop_WO_2
timestamp 1619646873
transform 1 0 1986 0 1 346
box -1 -64 165 57
use FlipFlop_WO  FlipFlop_WO_3
timestamp 1619646873
transform 1 0 1985 0 1 193
box -1 -64 165 57
use FlipFlop_WO  FlipFlop_WO_11
timestamp 1619646873
transform 0 -1 -99 1 0 -200
box -1 -64 165 57
use FlipFlop_WO  FlipFlop_WO_12
timestamp 1619646873
transform 0 -1 49 1 0 -200
box -1 -64 165 57
use FlipFlop_WO  FlipFlop_WO_4
timestamp 1619646873
transform 1 0 1984 0 1 21
box -1 -64 165 57
<< labels >>
rlabel metal2 -423 -68 -423 -68 3 a1
rlabel metal2 -423 -84 -423 -84 3 a2
rlabel metal2 -421 161 -421 161 1 a2
rlabel metal2 -425 462 -425 462 3 a3
rlabel metal2 -420 312 -420 312 1 b3
rlabel metal2 -421 613 -421 613 1 b4
rlabel metal2 -420 762 -420 762 1 a4
rlabel metal1 -428 537 -428 537 3 clk
rlabel metal2 330 -186 330 -186 1 vdd
rlabel metal2 526 -191 526 -191 1 gnd
rlabel space 2149 673 2149 673 7 Cout
rlabel space 2148 500 2148 500 7 s4
rlabel space 2149 338 2149 338 7 s3
rlabel space 2147 14 2147 14 7 s1
<< end >>
