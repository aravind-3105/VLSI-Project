* SPICE3 file created from 2NOR.ext - technology: scmos

.option scale=0.09u

M1000 a_13_5# B vdd w_0_n1# pfet w=40 l=2
+  ad=240 pd=92 as=200 ps=90
M1001 out A a_13_5# w_0_n1# pfet w=40 l=2
+  ad=280 pd=94 as=0 ps=0
M1002 out B gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=100 ps=60
M1003 gnd A out Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
C0 w_0_n1# gnd! 1.9fF
