* SPICE3 file created from CLA_With_FlipFlop.ext - technology: scmos

.option scale=0.09u

M1000 FlipFlop_WO_4/a_13_6# m1_1983_14# vdd FlipFlop_WO_4/w_0_0# pfet w=40 l=2
+  ad=240 pd=92 as=15860 ps=6926
M1001 FlipFlop_WO_4/a_13_n52# clk FlipFlop_WO_4/a_13_6# FlipFlop_WO_4/w_0_0# pfet w=40 l=2
+  ad=560 pd=108 as=0 ps=0
M1002 FlipFlop_WO_4/a_55_6# clk vdd FlipFlop_WO_4/w_0_0# pfet w=40 l=2
+  ad=680 pd=114 as=0 ps=0
M1003 FlipFlop_WO_4/a_90_6# FlipFlop_WO_4/a_55_6# vdd FlipFlop_WO_4/w_0_0# pfet w=40 l=2
+  ad=840 pd=202 as=0 ps=0
M1004 FlipFlop_WO_4/a_90_6# vdd vdd FlipFlop_WO_4/w_0_0# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 m1_2148_12# FlipFlop_WO_4/a_90_6# FlipFlop_WO_4/a_143_6# FlipFlop_WO_4/w_0_0# pfet w=40 l=2
+  ad=280 pd=94 as=280 ps=94
M1006 FlipFlop_WO_4/a_13_n52# m1_1983_14# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=9840 ps=4668
M1007 FlipFlop_WO_4/a_55_n52# clk gnd Gnd nfet w=20 l=2
+  ad=160 pd=56 as=0 ps=0
M1008 FlipFlop_WO_4/a_55_6# FlipFlop_WO_4/a_13_n52# FlipFlop_WO_4/a_55_n52# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1009 FlipFlop_WO_4/a_90_n52# FlipFlop_WO_4/a_55_6# gnd Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1010 FlipFlop_WO_4/a_90_6# FlipFlop_WO_4/a_94_n27# FlipFlop_WO_4/a_90_n52# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1011 m1_2148_12# FlipFlop_WO_4/a_90_6# gnd Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1012 FlipFlop_WO_12/a_13_6# FlipFlop_WO_12/a_9_n7# vdd FlipFlop_WO_12/w_0_0# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1013 FlipFlop_WO_12/a_13_n52# clk FlipFlop_WO_12/a_13_6# FlipFlop_WO_12/w_0_0# pfet w=40 l=2
+  ad=560 pd=108 as=0 ps=0
M1014 FlipFlop_WO_12/a_55_6# clk vdd FlipFlop_WO_12/w_0_0# pfet w=40 l=2
+  ad=680 pd=114 as=0 ps=0
M1015 FlipFlop_WO_12/a_90_6# FlipFlop_WO_12/a_55_6# vdd FlipFlop_WO_12/w_0_0# pfet w=40 l=2
+  ad=840 pd=202 as=0 ps=0
M1016 FlipFlop_WO_12/a_90_6# vdd vdd FlipFlop_WO_12/w_0_0# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1017 m1_n110_n21# FlipFlop_WO_12/a_90_6# FlipFlop_WO_12/a_143_6# FlipFlop_WO_12/w_0_0# pfet w=40 l=2
+  ad=280 pd=94 as=280 ps=94
M1018 FlipFlop_WO_12/a_13_n52# FlipFlop_WO_12/a_9_n7# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1019 FlipFlop_WO_12/a_55_n52# clk gnd Gnd nfet w=20 l=2
+  ad=160 pd=56 as=0 ps=0
M1020 FlipFlop_WO_12/a_55_6# FlipFlop_WO_12/a_13_n52# FlipFlop_WO_12/a_55_n52# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1021 FlipFlop_WO_12/a_90_n52# FlipFlop_WO_12/a_55_6# gnd Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1022 FlipFlop_WO_12/a_90_6# FlipFlop_WO_12/a_94_n27# FlipFlop_WO_12/a_90_n52# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1023 m1_n110_n21# FlipFlop_WO_12/a_90_6# gnd Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1024 FlipFlop_WO_11/a_13_6# a1 vdd FlipFlop_WO_11/w_0_0# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1025 FlipFlop_WO_11/a_13_n52# m1_n89_n203# FlipFlop_WO_11/a_13_6# FlipFlop_WO_11/w_0_0# pfet w=40 l=2
+  ad=560 pd=108 as=0 ps=0
M1026 FlipFlop_WO_11/a_55_6# m1_n89_n203# vdd FlipFlop_WO_11/w_0_0# pfet w=40 l=2
+  ad=680 pd=114 as=0 ps=0
M1027 FlipFlop_WO_11/a_90_6# FlipFlop_WO_11/a_55_6# vdd FlipFlop_WO_11/w_0_0# pfet w=40 l=2
+  ad=840 pd=202 as=0 ps=0
M1028 FlipFlop_WO_11/a_90_6# vdd vdd FlipFlop_WO_11/w_0_0# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1029 m2_n105_247# FlipFlop_WO_11/a_90_6# FlipFlop_WO_11/a_143_6# FlipFlop_WO_11/w_0_0# pfet w=40 l=2
+  ad=280 pd=94 as=280 ps=94
M1030 FlipFlop_WO_11/a_13_n52# a1 gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1031 FlipFlop_WO_11/a_55_n52# m1_n89_n203# gnd Gnd nfet w=20 l=2
+  ad=160 pd=56 as=0 ps=0
M1032 FlipFlop_WO_11/a_55_6# FlipFlop_WO_11/a_13_n52# FlipFlop_WO_11/a_55_n52# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1033 FlipFlop_WO_11/a_90_n52# FlipFlop_WO_11/a_55_6# gnd Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1034 FlipFlop_WO_11/a_90_6# FlipFlop_WO_11/a_94_n27# FlipFlop_WO_11/a_90_n52# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1035 m2_n105_247# FlipFlop_WO_11/a_90_6# gnd Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1036 FlipFlop_WO_3/a_13_6# m1_1978_186# vdd FlipFlop_WO_3/w_0_0# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1037 FlipFlop_WO_3/a_13_n52# clk FlipFlop_WO_3/a_13_6# FlipFlop_WO_3/w_0_0# pfet w=40 l=2
+  ad=560 pd=108 as=0 ps=0
M1038 FlipFlop_WO_3/a_55_6# clk vdd FlipFlop_WO_3/w_0_0# pfet w=40 l=2
+  ad=680 pd=114 as=0 ps=0
M1039 FlipFlop_WO_3/a_90_6# FlipFlop_WO_3/a_55_6# vdd FlipFlop_WO_3/w_0_0# pfet w=40 l=2
+  ad=840 pd=202 as=0 ps=0
M1040 FlipFlop_WO_3/a_90_6# vdd vdd FlipFlop_WO_3/w_0_0# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1041 FlipFlop_WO_3/a_152_n52# FlipFlop_WO_3/a_90_6# FlipFlop_WO_3/a_143_6# FlipFlop_WO_3/w_0_0# pfet w=40 l=2
+  ad=280 pd=94 as=280 ps=94
M1042 FlipFlop_WO_3/a_13_n52# m1_1978_186# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1043 FlipFlop_WO_3/a_55_n52# clk gnd Gnd nfet w=20 l=2
+  ad=160 pd=56 as=0 ps=0
M1044 FlipFlop_WO_3/a_55_6# FlipFlop_WO_3/a_13_n52# FlipFlop_WO_3/a_55_n52# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1045 FlipFlop_WO_3/a_90_n52# FlipFlop_WO_3/a_55_6# gnd Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1046 FlipFlop_WO_3/a_90_6# FlipFlop_WO_3/a_94_n27# FlipFlop_WO_3/a_90_n52# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1047 FlipFlop_WO_3/a_152_n52# FlipFlop_WO_3/a_90_6# gnd Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1048 FlipFlop_WO_2/a_13_6# m1_1978_339# vdd FlipFlop_WO_2/w_0_0# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1049 FlipFlop_WO_2/a_13_n52# clk FlipFlop_WO_2/a_13_6# FlipFlop_WO_2/w_0_0# pfet w=40 l=2
+  ad=560 pd=108 as=0 ps=0
M1050 FlipFlop_WO_2/a_55_6# clk vdd FlipFlop_WO_2/w_0_0# pfet w=40 l=2
+  ad=680 pd=114 as=0 ps=0
M1051 FlipFlop_WO_2/a_90_6# FlipFlop_WO_2/a_55_6# vdd FlipFlop_WO_2/w_0_0# pfet w=40 l=2
+  ad=840 pd=202 as=0 ps=0
M1052 FlipFlop_WO_2/a_90_6# vdd vdd FlipFlop_WO_2/w_0_0# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1053 m1_2150_337# FlipFlop_WO_2/a_90_6# FlipFlop_WO_2/a_143_6# FlipFlop_WO_2/w_0_0# pfet w=40 l=2
+  ad=280 pd=94 as=280 ps=94
M1054 FlipFlop_WO_2/a_13_n52# m1_1978_339# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1055 FlipFlop_WO_2/a_55_n52# clk gnd Gnd nfet w=20 l=2
+  ad=160 pd=56 as=0 ps=0
M1056 FlipFlop_WO_2/a_55_6# FlipFlop_WO_2/a_13_n52# FlipFlop_WO_2/a_55_n52# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1057 FlipFlop_WO_2/a_90_n52# FlipFlop_WO_2/a_55_6# gnd Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1058 FlipFlop_WO_2/a_90_6# FlipFlop_WO_2/a_94_n27# FlipFlop_WO_2/a_90_n52# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1059 m1_2150_337# FlipFlop_WO_2/a_90_6# gnd Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1060 FlipFlop_WO_1/a_13_6# m1_1939_499# vdd FlipFlop_WO_1/w_0_0# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1061 FlipFlop_WO_1/a_13_n52# clk FlipFlop_WO_1/a_13_6# FlipFlop_WO_1/w_0_0# pfet w=40 l=2
+  ad=560 pd=108 as=0 ps=0
M1062 FlipFlop_WO_1/a_55_6# clk vdd FlipFlop_WO_1/w_0_0# pfet w=40 l=2
+  ad=680 pd=114 as=0 ps=0
M1063 FlipFlop_WO_1/a_90_6# FlipFlop_WO_1/a_55_6# vdd FlipFlop_WO_1/w_0_0# pfet w=40 l=2
+  ad=840 pd=202 as=0 ps=0
M1064 FlipFlop_WO_1/a_90_6# vdd vdd FlipFlop_WO_1/w_0_0# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1065 m1_2149_498# FlipFlop_WO_1/a_90_6# FlipFlop_WO_1/a_143_6# FlipFlop_WO_1/w_0_0# pfet w=40 l=2
+  ad=280 pd=94 as=280 ps=94
M1066 FlipFlop_WO_1/a_13_n52# m1_1939_499# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1067 FlipFlop_WO_1/a_55_n52# clk gnd Gnd nfet w=20 l=2
+  ad=160 pd=56 as=0 ps=0
M1068 FlipFlop_WO_1/a_55_6# FlipFlop_WO_1/a_13_n52# FlipFlop_WO_1/a_55_n52# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1069 FlipFlop_WO_1/a_90_n52# FlipFlop_WO_1/a_55_6# gnd Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1070 FlipFlop_WO_1/a_90_6# FlipFlop_WO_1/a_94_n27# FlipFlop_WO_1/a_90_n52# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1071 m1_2149_498# FlipFlop_WO_1/a_90_6# gnd Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1072 FlipFlop_WO_0/a_13_6# m1_1015_205# vdd FlipFlop_WO_0/w_0_0# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1073 FlipFlop_WO_0/a_13_n52# clk FlipFlop_WO_0/a_13_6# FlipFlop_WO_0/w_0_0# pfet w=40 l=2
+  ad=560 pd=108 as=0 ps=0
M1074 FlipFlop_WO_0/a_55_6# clk vdd FlipFlop_WO_0/w_0_0# pfet w=40 l=2
+  ad=680 pd=114 as=0 ps=0
M1075 FlipFlop_WO_0/a_90_6# FlipFlop_WO_0/a_55_6# vdd FlipFlop_WO_0/w_0_0# pfet w=40 l=2
+  ad=840 pd=202 as=0 ps=0
M1076 FlipFlop_WO_0/a_90_6# vdd vdd FlipFlop_WO_0/w_0_0# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1077 m1_2150_671# FlipFlop_WO_0/a_90_6# FlipFlop_WO_0/a_143_6# FlipFlop_WO_0/w_0_0# pfet w=40 l=2
+  ad=280 pd=94 as=280 ps=94
M1078 FlipFlop_WO_0/a_13_n52# m1_1015_205# m1_1960_615# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=500 ps=210
M1079 FlipFlop_WO_0/a_55_n52# clk m1_1960_615# Gnd nfet w=20 l=2
+  ad=160 pd=56 as=0 ps=0
M1080 FlipFlop_WO_0/a_55_6# FlipFlop_WO_0/a_13_n52# FlipFlop_WO_0/a_55_n52# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1081 FlipFlop_WO_0/a_90_n52# FlipFlop_WO_0/a_55_6# m1_1960_615# Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1082 FlipFlop_WO_0/a_90_6# FlipFlop_WO_0/a_94_n27# FlipFlop_WO_0/a_90_n52# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1083 m1_2150_671# FlipFlop_WO_0/a_90_6# m1_1960_615# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1084 SUM_WO_0/XOR_WO_3/a_59_n30# m1_773_184# SUM_WO_0/XOR_WO_3/2INV_1/a_6_87# SUM_WO_0/XOR_WO_3/2INV_1/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1085 SUM_WO_0/XOR_WO_3/a_59_n30# m1_773_184# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1086 SUM_WO_0/XOR_WO_3/a_51_n59# m2_105_807# vdd SUM_WO_0/XOR_WO_3/2INV_0/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1087 SUM_WO_0/XOR_WO_3/a_51_n59# m2_105_807# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1088 vdd SUM_WO_0/XOR_WO_3/a_51_n59# SUM_WO_0/XOR_WO_3/a_56_27# SUM_WO_0/XOR_WO_3/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=400 ps=180
M1089 SUM_WO_0/XOR_WO_3/a_71_27# SUM_WO_0/XOR_WO_3/a_59_n30# vdd SUM_WO_0/XOR_WO_3/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1090 m1_1939_499# m2_105_807# SUM_WO_0/XOR_WO_3/a_71_27# SUM_WO_0/XOR_WO_3/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1091 SUM_WO_0/XOR_WO_3/a_56_27# m1_773_184# m1_1939_499# SUM_WO_0/XOR_WO_3/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1092 SUM_WO_0/XOR_WO_3/a_63_n51# SUM_WO_0/XOR_WO_3/a_59_n30# gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1093 m1_1939_499# SUM_WO_0/XOR_WO_3/a_51_n59# SUM_WO_0/XOR_WO_3/a_63_n51# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1094 SUM_WO_0/XOR_WO_3/a_79_n51# m2_105_807# m1_1939_499# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1095 gnd m1_773_184# SUM_WO_0/XOR_WO_3/a_79_n51# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1096 SUM_WO_0/XOR_WO_2/a_59_n30# m1_603_147# SUM_WO_0/XOR_WO_2/2INV_1/a_6_87# SUM_WO_0/XOR_WO_2/2INV_1/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1097 SUM_WO_0/XOR_WO_2/a_59_n30# m1_603_147# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1098 SUM_WO_0/XOR_WO_2/a_51_n59# m2_106_663# vdd SUM_WO_0/XOR_WO_2/2INV_0/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1099 SUM_WO_0/XOR_WO_2/a_51_n59# m2_106_663# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1100 vdd SUM_WO_0/XOR_WO_2/a_51_n59# SUM_WO_0/XOR_WO_2/a_56_27# SUM_WO_0/XOR_WO_2/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=400 ps=180
M1101 SUM_WO_0/XOR_WO_2/a_71_27# SUM_WO_0/XOR_WO_2/a_59_n30# vdd SUM_WO_0/XOR_WO_2/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1102 m1_1978_339# m2_106_663# SUM_WO_0/XOR_WO_2/a_71_27# SUM_WO_0/XOR_WO_2/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1103 SUM_WO_0/XOR_WO_2/a_56_27# m1_603_147# m1_1978_339# SUM_WO_0/XOR_WO_2/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1104 SUM_WO_0/XOR_WO_2/a_63_n51# SUM_WO_0/XOR_WO_2/a_59_n30# gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1105 m1_1978_339# SUM_WO_0/XOR_WO_2/a_51_n59# SUM_WO_0/XOR_WO_2/a_63_n51# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1106 SUM_WO_0/XOR_WO_2/a_79_n51# m2_106_663# m1_1978_339# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1107 gnd m1_603_147# SUM_WO_0/XOR_WO_2/a_79_n51# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1108 SUM_WO_0/XOR_WO_1/a_59_n30# m1_1395_46# SUM_WO_0/XOR_WO_1/2INV_1/a_6_87# SUM_WO_0/XOR_WO_1/2INV_1/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1109 SUM_WO_0/XOR_WO_1/a_59_n30# m1_1395_46# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1110 SUM_WO_0/XOR_WO_1/a_51_n59# m2_106_520# vdd SUM_WO_0/XOR_WO_1/2INV_0/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1111 SUM_WO_0/XOR_WO_1/a_51_n59# m2_106_520# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1112 vdd SUM_WO_0/XOR_WO_1/a_51_n59# SUM_WO_0/XOR_WO_1/a_56_27# SUM_WO_0/XOR_WO_1/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=400 ps=180
M1113 SUM_WO_0/XOR_WO_1/a_71_27# SUM_WO_0/XOR_WO_1/a_59_n30# vdd SUM_WO_0/XOR_WO_1/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1114 m1_1978_186# m2_106_520# SUM_WO_0/XOR_WO_1/a_71_27# SUM_WO_0/XOR_WO_1/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1115 SUM_WO_0/XOR_WO_1/a_56_27# m1_1395_46# m1_1978_186# SUM_WO_0/XOR_WO_1/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1116 SUM_WO_0/XOR_WO_1/a_63_n51# SUM_WO_0/XOR_WO_1/a_59_n30# gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1117 m1_1978_186# SUM_WO_0/XOR_WO_1/a_51_n59# SUM_WO_0/XOR_WO_1/a_63_n51# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1118 SUM_WO_0/XOR_WO_1/a_79_n51# m2_106_520# m1_1978_186# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1119 gnd m1_1395_46# SUM_WO_0/XOR_WO_1/a_79_n51# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1120 SUM_WO_0/XOR_WO_0/a_59_n30# gnd SUM_WO_0/XOR_WO_0/2INV_1/a_6_87# SUM_WO_0/XOR_WO_0/2INV_1/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1121 SUM_WO_0/XOR_WO_0/a_59_n30# gnd gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1122 SUM_WO_0/XOR_WO_0/a_51_n59# m2_189_369# vdd SUM_WO_0/XOR_WO_0/2INV_0/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1123 SUM_WO_0/XOR_WO_0/a_51_n59# m2_189_369# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1124 vdd SUM_WO_0/XOR_WO_0/a_51_n59# SUM_WO_0/XOR_WO_0/a_56_27# SUM_WO_0/XOR_WO_0/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=400 ps=180
M1125 SUM_WO_0/XOR_WO_0/a_71_27# SUM_WO_0/XOR_WO_0/a_59_n30# vdd SUM_WO_0/XOR_WO_0/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1126 m1_1983_14# m2_189_369# SUM_WO_0/XOR_WO_0/a_71_27# SUM_WO_0/XOR_WO_0/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1127 SUM_WO_0/XOR_WO_0/a_56_27# gnd m1_1983_14# SUM_WO_0/XOR_WO_0/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1128 SUM_WO_0/XOR_WO_0/a_63_n51# SUM_WO_0/XOR_WO_0/a_59_n30# gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1129 m1_1983_14# SUM_WO_0/XOR_WO_0/a_51_n59# SUM_WO_0/XOR_WO_0/a_63_n51# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1130 SUM_WO_0/XOR_WO_0/a_79_n51# m2_189_369# m1_1983_14# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1131 gnd gnd SUM_WO_0/XOR_WO_0/a_79_n51# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1132 m1_1015_205# Carry_WO_0/m1_409_n151# Carry_WO_0/2INV_8/a_6_87# Carry_WO_0/2INV_8/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1133 m1_1015_205# Carry_WO_0/m1_409_n151# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1134 Carry_WO_0/4NOR_WO_0/a_13_6# Carry_WO_0/m1_395_n85# vdd Carry_WO_0/4NOR_WO_0/w_0_0# pfet w=80 l=2
+  ad=480 pd=172 as=0 ps=0
M1135 Carry_WO_0/4NOR_WO_0/a_21_6# Carry_WO_0/m1_402_n83# Carry_WO_0/4NOR_WO_0/a_13_6# Carry_WO_0/4NOR_WO_0/w_0_0# pfet w=80 l=2
+  ad=480 pd=172 as=0 ps=0
M1136 Carry_WO_0/4NOR_WO_0/a_29_6# Carry_WO_0/m1_409_n82# Carry_WO_0/4NOR_WO_0/a_21_6# Carry_WO_0/4NOR_WO_0/w_0_0# pfet w=80 l=2
+  ad=480 pd=172 as=0 ps=0
M1137 Carry_WO_0/m1_409_n151# m1_243_38# Carry_WO_0/4NOR_WO_0/a_29_6# Carry_WO_0/4NOR_WO_0/w_0_0# pfet w=80 l=2
+  ad=560 pd=174 as=0 ps=0
M1138 Carry_WO_0/m1_409_n151# Carry_WO_0/m1_395_n85# gnd Gnd nfet w=10 l=2
+  ad=120 pd=64 as=0 ps=0
M1139 gnd Carry_WO_0/m1_402_n83# Carry_WO_0/m1_409_n151# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1140 Carry_WO_0/m1_409_n151# Carry_WO_0/m1_409_n82# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1141 gnd m1_243_38# Carry_WO_0/m1_409_n151# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1142 Carry_WO_0/m1_409_n82# Carry_WO_0/m1_683_20# Carry_WO_0/2INV_7/a_6_87# Carry_WO_0/2INV_7/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1143 Carry_WO_0/m1_409_n82# Carry_WO_0/m1_683_20# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1144 Carry_WO_0/m1_683_20# m2_105_807# vdd Carry_WO_0/4NAND_WO_0/w_0_0# pfet w=20 l=2
+  ad=240 pd=104 as=0 ps=0
M1145 vdd m2_106_663# Carry_WO_0/m1_683_20# Carry_WO_0/4NAND_WO_0/w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1146 Carry_WO_0/m1_683_20# m2_106_520# vdd Carry_WO_0/4NAND_WO_0/w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1147 vdd m1_1395_46# Carry_WO_0/m1_683_20# Carry_WO_0/4NAND_WO_0/w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1148 Carry_WO_0/4NAND_WO_0/a_13_n78# m2_105_807# gnd Gnd nfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1149 Carry_WO_0/4NAND_WO_0/a_21_n78# m2_106_663# Carry_WO_0/4NAND_WO_0/a_13_n78# Gnd nfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1150 Carry_WO_0/4NAND_WO_0/a_29_n78# m2_106_520# Carry_WO_0/4NAND_WO_0/a_21_n78# Gnd nfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1151 Carry_WO_0/m1_683_20# m1_1395_46# Carry_WO_0/4NAND_WO_0/a_29_n78# Gnd nfet w=40 l=2
+  ad=280 pd=94 as=0 ps=0
M1152 Carry_WO_0/3NOR_WO_0/a_14_3# Carry_WO_0/m1_174_23# vdd Carry_WO_0/3NOR_WO_0/w_1_n3# pfet w=60 l=2
+  ad=360 pd=132 as=0 ps=0
M1153 Carry_WO_0/3NOR_WO_0/a_22_3# m1_240_112# Carry_WO_0/3NOR_WO_0/a_14_3# Carry_WO_0/3NOR_WO_0/w_1_n3# pfet w=60 l=2
+  ad=360 pd=132 as=0 ps=0
M1154 Carry_WO_0/m1_194_n80# Carry_WO_0/m1_226_n94# Carry_WO_0/3NOR_WO_0/a_22_3# Carry_WO_0/3NOR_WO_0/w_1_n3# pfet w=60 l=2
+  ad=420 pd=134 as=0 ps=0
M1155 Carry_WO_0/m1_194_n80# Carry_WO_0/m1_174_23# gnd Gnd nfet w=10 l=2
+  ad=130 pd=66 as=0 ps=0
M1156 gnd m1_240_112# Carry_WO_0/m1_194_n80# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1157 Carry_WO_0/m1_194_n80# Carry_WO_0/m1_226_n94# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1158 m1_773_184# Carry_WO_0/m1_194_n80# Carry_WO_0/2INV_3/a_6_87# Carry_WO_0/2INV_3/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1159 m1_773_184# Carry_WO_0/m1_194_n80# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1160 Carry_WO_0/m1_402_n83# Carry_WO_0/m1_526_53# Carry_WO_0/2INV_6/a_6_87# Carry_WO_0/2INV_6/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1161 Carry_WO_0/m1_402_n83# Carry_WO_0/m1_526_53# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1162 Carry_WO_0/m1_526_53# m2_105_807# vdd Carry_WO_0/3NAND_WO_1/w_0_0# pfet w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M1163 vdd m2_106_663# Carry_WO_0/m1_526_53# Carry_WO_0/3NAND_WO_1/w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1164 Carry_WO_0/m1_526_53# m1_240_299# vdd Carry_WO_0/3NAND_WO_1/w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1165 Carry_WO_0/3NAND_WO_1/a_13_n61# m2_105_807# gnd Gnd nfet w=30 l=2
+  ad=180 pd=72 as=0 ps=0
M1166 Carry_WO_0/3NAND_WO_1/a_21_n61# m2_106_663# Carry_WO_0/3NAND_WO_1/a_13_n61# Gnd nfet w=30 l=2
+  ad=180 pd=72 as=0 ps=0
M1167 Carry_WO_0/m1_526_53# m1_240_299# Carry_WO_0/3NAND_WO_1/a_21_n61# Gnd nfet w=30 l=2
+  ad=210 pd=74 as=0 ps=0
M1168 Carry_WO_0/m1_395_n85# Carry_WO_0/m1_398_36# Carry_WO_0/2INV_5/a_6_87# Carry_WO_0/2INV_5/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1169 Carry_WO_0/m1_395_n85# Carry_WO_0/m1_398_36# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1170 Carry_WO_0/m1_398_36# m2_105_807# vdd Carry_WO_0/2NAND_WO_2/w_0_0# pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1171 vdd m1_240_112# Carry_WO_0/m1_398_36# Carry_WO_0/2NAND_WO_2/w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1172 Carry_WO_0/2NAND_WO_2/a_13_n43# m2_105_807# gnd Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1173 Carry_WO_0/m1_398_36# m1_240_112# Carry_WO_0/2NAND_WO_2/a_13_n43# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1174 Carry_WO_0/m1_226_n94# Carry_WO_0/m1_252_46# Carry_WO_0/2INV_4/a_6_87# Carry_WO_0/2INV_4/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1175 Carry_WO_0/m1_226_n94# Carry_WO_0/m1_252_46# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1176 Carry_WO_0/m1_252_46# m1_1395_46# vdd Carry_WO_0/3NAND_WO_0/w_0_0# pfet w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M1177 vdd m2_106_520# Carry_WO_0/m1_252_46# Carry_WO_0/3NAND_WO_0/w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1178 Carry_WO_0/m1_252_46# m2_106_663# vdd Carry_WO_0/3NAND_WO_0/w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1179 Carry_WO_0/3NAND_WO_0/a_13_n61# m1_1395_46# gnd Gnd nfet w=30 l=2
+  ad=180 pd=72 as=0 ps=0
M1180 Carry_WO_0/3NAND_WO_0/a_21_n61# m2_106_520# Carry_WO_0/3NAND_WO_0/a_13_n61# Gnd nfet w=30 l=2
+  ad=180 pd=72 as=0 ps=0
M1181 Carry_WO_0/m1_252_46# m2_106_663# Carry_WO_0/3NAND_WO_0/a_21_n61# Gnd nfet w=30 l=2
+  ad=210 pd=74 as=0 ps=0
M1182 Carry_WO_0/m1_174_23# Carry_WO_0/m1_145_29# Carry_WO_0/2INV_2/a_6_87# Carry_WO_0/2INV_2/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1183 Carry_WO_0/m1_174_23# Carry_WO_0/m1_145_29# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1184 Carry_WO_0/m1_145_29# m2_106_663# vdd Carry_WO_0/2NAND_WO_1/w_0_0# pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1185 vdd m1_240_299# Carry_WO_0/m1_145_29# Carry_WO_0/2NAND_WO_1/w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1186 Carry_WO_0/2NAND_WO_1/a_13_n43# m2_106_663# gnd Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1187 Carry_WO_0/m1_145_29# m1_240_299# Carry_WO_0/2NAND_WO_1/a_13_n43# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1188 Carry_WO_0/2NOR_WO_0/a_13_5# Carry_WO_0/m1_63_n31# vdd Carry_WO_0/w_38_n91# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1189 Carry_WO_0/m1_19_n37# m1_240_299# Carry_WO_0/2NOR_WO_0/a_13_5# Carry_WO_0/w_38_n91# pfet w=40 l=2
+  ad=280 pd=94 as=0 ps=0
M1190 Carry_WO_0/m1_19_n37# Carry_WO_0/m1_63_n31# gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1191 gnd m1_240_299# Carry_WO_0/m1_19_n37# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1192 m1_603_147# Carry_WO_0/m1_19_n37# Carry_WO_0/2INV_1/a_6_87# Carry_WO_0/2INV_1/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1193 m1_603_147# Carry_WO_0/m1_19_n37# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1194 Carry_WO_0/m1_63_n31# Carry_WO_0/m1_25_30# Carry_WO_0/2INV_0/a_6_87# Carry_WO_0/2INV_0/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1195 Carry_WO_0/m1_63_n31# Carry_WO_0/m1_25_30# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1196 Carry_WO_0/m1_25_30# m1_1395_46# vdd Carry_WO_0/w_7_77# pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1197 vdd m2_106_520# Carry_WO_0/m1_25_30# Carry_WO_0/w_7_77# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1198 Carry_WO_0/2NAND_WO_0/a_13_n43# m1_1395_46# gnd Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1199 Carry_WO_0/m1_25_30# m2_106_520# Carry_WO_0/2NAND_WO_0/a_13_n43# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1200 m1_240_299# m1_195_305# PropagateGenerate_WO_0/2INV_3/a_6_87# PropagateGenerate_WO_0/2INV_3/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1201 m1_240_299# m1_195_305# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1202 m1_1395_46# m1_201_222# PropagateGenerate_WO_0/2INV_2/a_6_87# PropagateGenerate_WO_0/2INV_2/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1203 m1_1395_46# m1_201_222# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1204 m1_240_112# m1_199_103# PropagateGenerate_WO_0/2INV_1/a_6_87# PropagateGenerate_WO_0/2INV_1/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1205 m1_240_112# m1_199_103# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1206 m1_243_38# m1_195_44# PropagateGenerate_WO_0/2INV_0/a_6_87# PropagateGenerate_WO_0/2INV_0/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1207 m1_243_38# m1_195_44# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1208 PropagateGenerate_WO_0/XOR_WO_3/a_59_n30# m1_n185_609# PropagateGenerate_WO_0/XOR_WO_3/2INV_1/a_6_87# PropagateGenerate_WO_0/XOR_WO_3/2INV_1/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1209 PropagateGenerate_WO_0/XOR_WO_3/a_59_n30# m1_n185_609# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1210 PropagateGenerate_WO_0/XOR_WO_3/a_51_n59# m1_n188_758# vdd PropagateGenerate_WO_0/XOR_WO_3/2INV_0/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1211 PropagateGenerate_WO_0/XOR_WO_3/a_51_n59# m1_n188_758# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1212 vdd PropagateGenerate_WO_0/XOR_WO_3/a_51_n59# PropagateGenerate_WO_0/XOR_WO_3/a_56_27# PropagateGenerate_WO_0/XOR_WO_3/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=400 ps=180
M1213 PropagateGenerate_WO_0/XOR_WO_3/a_71_27# PropagateGenerate_WO_0/XOR_WO_3/a_59_n30# vdd PropagateGenerate_WO_0/XOR_WO_3/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1214 m2_105_807# m1_n188_758# PropagateGenerate_WO_0/XOR_WO_3/a_71_27# PropagateGenerate_WO_0/XOR_WO_3/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1215 PropagateGenerate_WO_0/XOR_WO_3/a_56_27# m1_n185_609# m2_105_807# PropagateGenerate_WO_0/XOR_WO_3/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1216 PropagateGenerate_WO_0/XOR_WO_3/a_63_n51# PropagateGenerate_WO_0/XOR_WO_3/a_59_n30# gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1217 m2_105_807# PropagateGenerate_WO_0/XOR_WO_3/a_51_n59# PropagateGenerate_WO_0/XOR_WO_3/a_63_n51# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1218 PropagateGenerate_WO_0/XOR_WO_3/a_79_n51# m1_n188_758# m2_105_807# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1219 gnd m1_n185_609# PropagateGenerate_WO_0/XOR_WO_3/a_79_n51# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1220 PropagateGenerate_WO_0/XOR_WO_2/a_59_n30# m1_n188_308# PropagateGenerate_WO_0/XOR_WO_2/2INV_1/a_6_87# PropagateGenerate_WO_0/XOR_WO_2/2INV_1/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1221 PropagateGenerate_WO_0/XOR_WO_2/a_59_n30# m1_n188_308# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1222 PropagateGenerate_WO_0/XOR_WO_2/a_51_n59# m1_n193_459# vdd PropagateGenerate_WO_0/XOR_WO_2/2INV_0/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1223 PropagateGenerate_WO_0/XOR_WO_2/a_51_n59# m1_n193_459# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1224 vdd PropagateGenerate_WO_0/XOR_WO_2/a_51_n59# PropagateGenerate_WO_0/XOR_WO_2/a_56_27# PropagateGenerate_WO_0/XOR_WO_2/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=400 ps=180
M1225 PropagateGenerate_WO_0/XOR_WO_2/a_71_27# PropagateGenerate_WO_0/XOR_WO_2/a_59_n30# vdd PropagateGenerate_WO_0/XOR_WO_2/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1226 m2_106_663# m1_n193_459# PropagateGenerate_WO_0/XOR_WO_2/a_71_27# PropagateGenerate_WO_0/XOR_WO_2/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1227 PropagateGenerate_WO_0/XOR_WO_2/a_56_27# m1_n188_308# m2_106_663# PropagateGenerate_WO_0/XOR_WO_2/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1228 PropagateGenerate_WO_0/XOR_WO_2/a_63_n51# PropagateGenerate_WO_0/XOR_WO_2/a_59_n30# gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1229 m2_106_663# PropagateGenerate_WO_0/XOR_WO_2/a_51_n59# PropagateGenerate_WO_0/XOR_WO_2/a_63_n51# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1230 PropagateGenerate_WO_0/XOR_WO_2/a_79_n51# m1_n193_459# m2_106_663# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1231 gnd m1_n188_308# PropagateGenerate_WO_0/XOR_WO_2/a_79_n51# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1232 PropagateGenerate_WO_0/XOR_WO_1/a_59_n30# m1_n188_6# PropagateGenerate_WO_0/XOR_WO_1/2INV_1/a_6_87# PropagateGenerate_WO_0/XOR_WO_1/2INV_1/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1233 PropagateGenerate_WO_0/XOR_WO_1/a_59_n30# m1_n188_6# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1234 PropagateGenerate_WO_0/XOR_WO_1/a_51_n59# m2_n89_397# vdd PropagateGenerate_WO_0/XOR_WO_1/2INV_0/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1235 PropagateGenerate_WO_0/XOR_WO_1/a_51_n59# m2_n89_397# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1236 vdd PropagateGenerate_WO_0/XOR_WO_1/a_51_n59# PropagateGenerate_WO_0/XOR_WO_1/a_56_27# PropagateGenerate_WO_0/XOR_WO_1/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=400 ps=180
M1237 PropagateGenerate_WO_0/XOR_WO_1/a_71_27# PropagateGenerate_WO_0/XOR_WO_1/a_59_n30# vdd PropagateGenerate_WO_0/XOR_WO_1/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1238 m2_106_520# m2_n89_397# PropagateGenerate_WO_0/XOR_WO_1/a_71_27# PropagateGenerate_WO_0/XOR_WO_1/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1239 PropagateGenerate_WO_0/XOR_WO_1/a_56_27# m1_n188_6# m2_106_520# PropagateGenerate_WO_0/XOR_WO_1/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1240 PropagateGenerate_WO_0/XOR_WO_1/a_63_n51# PropagateGenerate_WO_0/XOR_WO_1/a_59_n30# gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1241 m2_106_520# PropagateGenerate_WO_0/XOR_WO_1/a_51_n59# PropagateGenerate_WO_0/XOR_WO_1/a_63_n51# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1242 PropagateGenerate_WO_0/XOR_WO_1/a_79_n51# m2_n89_397# m2_106_520# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1243 gnd m1_n188_6# PropagateGenerate_WO_0/XOR_WO_1/a_79_n51# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1244 PropagateGenerate_WO_0/XOR_WO_0/a_59_n30# m1_n110_n21# PropagateGenerate_WO_0/XOR_WO_0/2INV_1/a_6_87# PropagateGenerate_WO_0/XOR_WO_0/2INV_1/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1245 PropagateGenerate_WO_0/XOR_WO_0/a_59_n30# m1_n110_n21# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1246 PropagateGenerate_WO_0/XOR_WO_0/a_51_n59# m2_n105_247# vdd PropagateGenerate_WO_0/XOR_WO_0/2INV_0/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1247 PropagateGenerate_WO_0/XOR_WO_0/a_51_n59# m2_n105_247# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1248 vdd PropagateGenerate_WO_0/XOR_WO_0/a_51_n59# PropagateGenerate_WO_0/XOR_WO_0/a_56_27# PropagateGenerate_WO_0/XOR_WO_0/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=400 ps=180
M1249 PropagateGenerate_WO_0/XOR_WO_0/a_71_27# PropagateGenerate_WO_0/XOR_WO_0/a_59_n30# vdd PropagateGenerate_WO_0/XOR_WO_0/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1250 m2_189_369# m2_n105_247# PropagateGenerate_WO_0/XOR_WO_0/a_71_27# PropagateGenerate_WO_0/XOR_WO_0/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1251 PropagateGenerate_WO_0/XOR_WO_0/a_56_27# m1_n110_n21# m2_189_369# PropagateGenerate_WO_0/XOR_WO_0/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1252 PropagateGenerate_WO_0/XOR_WO_0/a_63_n51# PropagateGenerate_WO_0/XOR_WO_0/a_59_n30# gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1253 m2_189_369# PropagateGenerate_WO_0/XOR_WO_0/a_51_n59# PropagateGenerate_WO_0/XOR_WO_0/a_63_n51# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1254 PropagateGenerate_WO_0/XOR_WO_0/a_79_n51# m2_n105_247# m2_189_369# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1255 gnd m1_n110_n21# PropagateGenerate_WO_0/XOR_WO_0/a_79_n51# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1256 m1_195_305# m2_n89_397# vdd PropagateGenerate_WO_0/2AND_WO_1/w_0_0# pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1257 vdd m1_n188_6# m1_195_305# PropagateGenerate_WO_0/2AND_WO_1/w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1258 PropagateGenerate_WO_0/2AND_WO_1/a_13_n43# m2_n89_397# gnd Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1259 m1_195_305# m1_n188_6# PropagateGenerate_WO_0/2AND_WO_1/a_13_n43# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1260 m1_195_44# m1_n188_758# vdd PropagateGenerate_WO_0/2AND_WO_3/w_0_0# pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1261 vdd m1_n185_609# m1_195_44# PropagateGenerate_WO_0/2AND_WO_3/w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1262 PropagateGenerate_WO_0/2AND_WO_3/a_13_n43# m1_n188_758# gnd Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1263 m1_195_44# m1_n185_609# PropagateGenerate_WO_0/2AND_WO_3/a_13_n43# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1264 m1_201_222# m2_n105_247# vdd PropagateGenerate_WO_0/2AND_WO_0/w_0_0# pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1265 vdd m1_n110_n21# m1_201_222# PropagateGenerate_WO_0/2AND_WO_0/w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1266 PropagateGenerate_WO_0/2AND_WO_0/a_13_n43# m2_n105_247# gnd Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1267 m1_201_222# m1_n110_n21# PropagateGenerate_WO_0/2AND_WO_0/a_13_n43# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1268 m1_199_103# m1_n193_459# vdd PropagateGenerate_WO_0/2AND_WO_2/w_0_0# pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1269 vdd m1_n188_308# m1_199_103# PropagateGenerate_WO_0/2AND_WO_2/w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1270 PropagateGenerate_WO_0/2AND_WO_2/a_13_n43# m1_n193_459# gnd Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1271 m1_199_103# m1_n188_308# PropagateGenerate_WO_0/2AND_WO_2/a_13_n43# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1272 FlipFlop_WO_10/a_13_6# m1_n353_8# vdd FlipFlop_WO_10/w_0_0# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1273 FlipFlop_WO_10/a_13_n52# clk FlipFlop_WO_10/a_13_6# FlipFlop_WO_10/w_0_0# pfet w=40 l=2
+  ad=560 pd=108 as=0 ps=0
M1274 FlipFlop_WO_10/a_55_6# clk vdd FlipFlop_WO_10/w_0_0# pfet w=40 l=2
+  ad=680 pd=114 as=0 ps=0
M1275 FlipFlop_WO_10/a_90_6# FlipFlop_WO_10/a_55_6# vdd FlipFlop_WO_10/w_0_0# pfet w=40 l=2
+  ad=840 pd=202 as=0 ps=0
M1276 FlipFlop_WO_10/a_90_6# vdd vdd FlipFlop_WO_10/w_0_0# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1277 m1_n188_6# FlipFlop_WO_10/a_90_6# FlipFlop_WO_10/a_143_6# FlipFlop_WO_10/w_0_0# pfet w=40 l=2
+  ad=280 pd=94 as=280 ps=94
M1278 FlipFlop_WO_10/a_13_n52# m1_n353_8# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1279 FlipFlop_WO_10/a_55_n52# clk gnd Gnd nfet w=20 l=2
+  ad=160 pd=56 as=0 ps=0
M1280 FlipFlop_WO_10/a_55_6# FlipFlop_WO_10/a_13_n52# FlipFlop_WO_10/a_55_n52# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1281 FlipFlop_WO_10/a_90_n52# FlipFlop_WO_10/a_55_6# gnd Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1282 FlipFlop_WO_10/a_90_6# FlipFlop_WO_10/a_94_n27# FlipFlop_WO_10/a_90_n52# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1283 m1_n188_6# FlipFlop_WO_10/a_90_6# gnd Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1284 FlipFlop_WO_9/a_13_6# a2 vdd FlipFlop_WO_9/w_0_0# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1285 FlipFlop_WO_9/a_13_n52# clk FlipFlop_WO_9/a_13_6# FlipFlop_WO_9/w_0_0# pfet w=40 l=2
+  ad=560 pd=108 as=0 ps=0
M1286 FlipFlop_WO_9/a_55_6# clk vdd FlipFlop_WO_9/w_0_0# pfet w=40 l=2
+  ad=680 pd=114 as=0 ps=0
M1287 FlipFlop_WO_9/a_90_6# FlipFlop_WO_9/a_55_6# vdd FlipFlop_WO_9/w_0_0# pfet w=40 l=2
+  ad=840 pd=202 as=0 ps=0
M1288 FlipFlop_WO_9/a_90_6# vdd vdd FlipFlop_WO_9/w_0_0# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1289 m2_n89_397# FlipFlop_WO_9/a_90_6# FlipFlop_WO_9/a_143_6# FlipFlop_WO_9/w_0_0# pfet w=40 l=2
+  ad=280 pd=94 as=280 ps=94
M1290 FlipFlop_WO_9/a_13_n52# a2 gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1291 FlipFlop_WO_9/a_55_n52# clk gnd Gnd nfet w=20 l=2
+  ad=160 pd=56 as=0 ps=0
M1292 FlipFlop_WO_9/a_55_6# FlipFlop_WO_9/a_13_n52# FlipFlop_WO_9/a_55_n52# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1293 FlipFlop_WO_9/a_90_n52# FlipFlop_WO_9/a_55_6# gnd Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1294 FlipFlop_WO_9/a_90_6# FlipFlop_WO_9/a_94_n27# FlipFlop_WO_9/a_90_n52# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1295 m2_n89_397# FlipFlop_WO_9/a_90_6# gnd Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1296 FlipFlop_WO_8/a_13_6# b3 FlipFlop_WO_8/a_6_6# FlipFlop_WO_8/w_0_0# pfet w=40 l=2
+  ad=240 pd=92 as=840 ps=362
M1297 FlipFlop_WO_8/a_13_n52# clk FlipFlop_WO_8/a_13_6# FlipFlop_WO_8/w_0_0# pfet w=40 l=2
+  ad=560 pd=108 as=0 ps=0
M1298 FlipFlop_WO_8/a_55_6# clk FlipFlop_WO_8/a_6_6# FlipFlop_WO_8/w_0_0# pfet w=40 l=2
+  ad=680 pd=114 as=0 ps=0
M1299 FlipFlop_WO_8/a_90_6# FlipFlop_WO_8/a_55_6# FlipFlop_WO_8/a_6_6# FlipFlop_WO_8/w_0_0# pfet w=40 l=2
+  ad=840 pd=202 as=0 ps=0
M1300 FlipFlop_WO_8/a_90_6# FlipFlop_WO_8/a_6_6# FlipFlop_WO_8/a_6_6# FlipFlop_WO_8/w_0_0# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1301 m1_n188_308# FlipFlop_WO_8/a_90_6# FlipFlop_WO_8/a_143_6# FlipFlop_WO_8/w_0_0# pfet w=40 l=2
+  ad=280 pd=94 as=280 ps=94
M1302 FlipFlop_WO_8/a_13_n52# b3 gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1303 FlipFlop_WO_8/a_55_n52# clk gnd Gnd nfet w=20 l=2
+  ad=160 pd=56 as=0 ps=0
M1304 FlipFlop_WO_8/a_55_6# FlipFlop_WO_8/a_13_n52# FlipFlop_WO_8/a_55_n52# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1305 FlipFlop_WO_8/a_90_n52# FlipFlop_WO_8/a_55_6# gnd Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1306 FlipFlop_WO_8/a_90_6# FlipFlop_WO_8/a_94_n27# FlipFlop_WO_8/a_90_n52# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1307 m1_n188_308# FlipFlop_WO_8/a_90_6# gnd Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1308 FlipFlop_WO_7/a_13_6# a3 vdd FlipFlop_WO_7/w_0_0# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1309 FlipFlop_WO_7/a_13_n52# clk FlipFlop_WO_7/a_13_6# FlipFlop_WO_7/w_0_0# pfet w=40 l=2
+  ad=560 pd=108 as=0 ps=0
M1310 FlipFlop_WO_7/a_55_6# clk vdd FlipFlop_WO_7/w_0_0# pfet w=40 l=2
+  ad=680 pd=114 as=0 ps=0
M1311 FlipFlop_WO_7/a_90_6# FlipFlop_WO_7/a_55_6# vdd FlipFlop_WO_7/w_0_0# pfet w=40 l=2
+  ad=840 pd=202 as=0 ps=0
M1312 FlipFlop_WO_7/a_90_6# vdd vdd FlipFlop_WO_7/w_0_0# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1313 m1_n193_459# FlipFlop_WO_7/a_90_6# FlipFlop_WO_7/a_143_6# FlipFlop_WO_7/w_0_0# pfet w=40 l=2
+  ad=280 pd=94 as=280 ps=94
M1314 FlipFlop_WO_7/a_13_n52# a3 gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1315 FlipFlop_WO_7/a_55_n52# clk gnd Gnd nfet w=20 l=2
+  ad=160 pd=56 as=0 ps=0
M1316 FlipFlop_WO_7/a_55_6# FlipFlop_WO_7/a_13_n52# FlipFlop_WO_7/a_55_n52# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1317 FlipFlop_WO_7/a_90_n52# FlipFlop_WO_7/a_55_6# gnd Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1318 FlipFlop_WO_7/a_90_6# FlipFlop_WO_7/a_94_n27# FlipFlop_WO_7/a_90_n52# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1319 m1_n193_459# FlipFlop_WO_7/a_90_6# gnd Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1320 FlipFlop_WO_6/a_13_6# b4 vdd FlipFlop_WO_6/w_0_0# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1321 FlipFlop_WO_6/a_13_n52# clk FlipFlop_WO_6/a_13_6# FlipFlop_WO_6/w_0_0# pfet w=40 l=2
+  ad=560 pd=108 as=0 ps=0
M1322 FlipFlop_WO_6/a_55_6# clk vdd FlipFlop_WO_6/w_0_0# pfet w=40 l=2
+  ad=680 pd=114 as=0 ps=0
M1323 FlipFlop_WO_6/a_90_6# FlipFlop_WO_6/a_55_6# vdd FlipFlop_WO_6/w_0_0# pfet w=40 l=2
+  ad=840 pd=202 as=0 ps=0
M1324 FlipFlop_WO_6/a_90_6# vdd vdd FlipFlop_WO_6/w_0_0# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1325 m1_n185_609# FlipFlop_WO_6/a_90_6# FlipFlop_WO_6/a_143_6# FlipFlop_WO_6/w_0_0# pfet w=40 l=2
+  ad=280 pd=94 as=280 ps=94
M1326 FlipFlop_WO_6/a_13_n52# b4 gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1327 FlipFlop_WO_6/a_55_n52# clk gnd Gnd nfet w=20 l=2
+  ad=160 pd=56 as=0 ps=0
M1328 FlipFlop_WO_6/a_55_6# FlipFlop_WO_6/a_13_n52# FlipFlop_WO_6/a_55_n52# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1329 FlipFlop_WO_6/a_90_n52# FlipFlop_WO_6/a_55_6# gnd Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1330 FlipFlop_WO_6/a_90_6# FlipFlop_WO_6/a_94_n27# FlipFlop_WO_6/a_90_n52# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1331 m1_n185_609# FlipFlop_WO_6/a_90_6# gnd Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1332 FlipFlop_WO_5/a_13_6# a4 vdd FlipFlop_WO_5/w_0_0# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1333 FlipFlop_WO_5/a_13_n52# clk FlipFlop_WO_5/a_13_6# FlipFlop_WO_5/w_0_0# pfet w=40 l=2
+  ad=560 pd=108 as=0 ps=0
M1334 FlipFlop_WO_5/a_55_6# clk vdd FlipFlop_WO_5/w_0_0# pfet w=40 l=2
+  ad=680 pd=114 as=0 ps=0
M1335 FlipFlop_WO_5/a_90_6# FlipFlop_WO_5/a_55_6# vdd FlipFlop_WO_5/w_0_0# pfet w=40 l=2
+  ad=840 pd=202 as=0 ps=0
M1336 FlipFlop_WO_5/a_90_6# vdd vdd FlipFlop_WO_5/w_0_0# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1337 m1_n188_758# FlipFlop_WO_5/a_90_6# FlipFlop_WO_5/a_143_6# FlipFlop_WO_5/w_0_0# pfet w=40 l=2
+  ad=280 pd=94 as=280 ps=94
M1338 FlipFlop_WO_5/a_13_n52# a4 gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1339 FlipFlop_WO_5/a_55_n52# clk gnd Gnd nfet w=20 l=2
+  ad=160 pd=56 as=0 ps=0
M1340 FlipFlop_WO_5/a_55_6# FlipFlop_WO_5/a_13_n52# FlipFlop_WO_5/a_55_n52# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1341 FlipFlop_WO_5/a_90_n52# FlipFlop_WO_5/a_55_6# gnd Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1342 FlipFlop_WO_5/a_90_6# FlipFlop_WO_5/a_94_n27# FlipFlop_WO_5/a_90_n52# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1343 m1_n188_758# FlipFlop_WO_5/a_90_6# gnd Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
C0 vdd m1_1395_46# 1.3fF
C1 FlipFlop_WO_8/w_0_0# FlipFlop_WO_8/a_6_6# 1.3fF
C2 SUM_WO_0/XOR_WO_3/a_56_27# m1_1939_499# 1.1fF
C3 m2_106_520# m2_106_663# 4.7fF
C4 m2_106_520# PropagateGenerate_WO_0/XOR_WO_1/a_56_27# 1.1fF
C5 SUM_WO_0/XOR_WO_0/a_56_27# m1_1983_14# 1.1fF
C6 FlipFlop_WO_4/w_0_0# vdd 1.3fF
C7 vdd m1_201_222# 1.2fF
C8 m2_105_807# PropagateGenerate_WO_0/XOR_WO_3/a_56_27# 1.1fF
C9 SUM_WO_0/XOR_WO_2/a_56_27# m1_1978_339# 1.1fF
C10 m1_240_299# m2_106_663# 6.4fF
C11 FlipFlop_WO_2/w_0_0# vdd 1.3fF
C12 Carry_WO_0/m1_402_n83# Carry_WO_0/m1_395_n85# 1.5fF
C13 vdd FlipFlop_WO_6/w_0_0# 1.3fF
C14 clk gnd 1.3fF
C15 Carry_WO_0/m1_409_n82# Carry_WO_0/m1_402_n83# 2.3fF
C16 PropagateGenerate_WO_0/XOR_WO_0/a_56_27# m2_189_369# 1.1fF
C17 vdd FlipFlop_WO_7/w_0_0# 1.3fF
C18 m2_189_369# gnd 2.3fF
C19 vdd FlipFlop_WO_10/w_0_0# 1.3fF
C20 m1_n185_609# m1_n188_758# 12.7fF
C21 m1_n193_459# m1_n188_308# 8.6fF
C22 FlipFlop_WO_12/w_0_0# vdd 1.3fF
C23 m2_106_520# m1_240_299# 2.5fF
C24 m1_1015_205# clk 1.1fF
C25 vdd m2_106_663# 1.1fF
C26 m2_106_520# m1_1395_46# 10.3fF
C27 m1_773_184# m2_105_807# 2.0fF
C28 vdd FlipFlop_WO_9/w_0_0# 1.3fF
C29 m2_105_807# m2_106_663# 4.3fF
C30 vdd gnd 2.1fF
C31 m1_240_112# Carry_WO_0/m1_226_n94# 1.1fF
C32 m1_240_112# m2_105_807# 2.9fF
C33 FlipFlop_WO_0/w_0_0# vdd 1.3fF
C34 m1_243_38# m2_105_807# 2.0fF
C35 m2_n105_247# m1_n110_n21# 3.7fF
C36 vdd FlipFlop_WO_5/w_0_0# 1.3fF
C37 vdd m1_n110_n21# 1.3fF
C38 m1_240_112# m2_106_663# 2.1fF
C39 FlipFlop_WO_3/w_0_0# vdd 1.3fF
C40 m2_n89_397# m1_n188_6# 6.1fF
C41 FlipFlop_WO_1/w_0_0# vdd 1.3fF
C42 m1_1015_205# vdd 2.1fF
C43 m1_243_38# m1_240_112# 2.0fF
C44 PropagateGenerate_WO_0/XOR_WO_2/a_56_27# m2_106_663# 1.1fF
C45 m1_n193_459# m1_n188_6# 2.4fF
C46 m1_240_299# Carry_WO_0/m1_63_n31# 1.2fF
C47 FlipFlop_WO_11/w_0_0# vdd 1.3fF
C48 m1_603_147# m2_106_663# 2.0fF
C49 m1_n188_308# m1_n188_758# 5.2fF
C50 SUM_WO_0/XOR_WO_1/a_56_27# m1_1978_186# 1.1fF
C51 m1_243_38# Carry_WO_0/m1_409_n82# 2.9fF
C52 gnd gnd! 85.0fF
C53 m1_n188_758# gnd! 7.1fF
C54 clk gnd! 32.4fF
C55 a4 gnd! 1.0fF
C56 FlipFlop_WO_5/w_0_0# gnd! 9.4fF
C57 b4 gnd! 1.1fF
C58 FlipFlop_WO_6/w_0_0# gnd! 9.4fF
C59 a3 gnd! 1.1fF
C60 FlipFlop_WO_7/w_0_0# gnd! 9.4fF
C61 b3 gnd! 1.1fF
C62 FlipFlop_WO_8/w_0_0# gnd! 9.4fF
C63 a2 gnd! 8.1fF
C64 FlipFlop_WO_9/w_0_0# gnd! 9.4fF
C65 m1_n353_8# gnd! 1.0fF
C66 FlipFlop_WO_10/w_0_0# gnd! 9.4fF
C67 m1_199_103# gnd! 1.4fF
C68 m1_n188_308# gnd! 6.6fF
C69 PropagateGenerate_WO_0/2AND_WO_2/w_0_0# gnd! 1.0fF
C70 m1_201_222# gnd! 1.1fF
C71 m1_n110_n21# gnd! 5.6fF
C72 PropagateGenerate_WO_0/2AND_WO_0/w_0_0# gnd! 1.0fF
C73 m1_n185_609# gnd! 7.9fF
C74 PropagateGenerate_WO_0/2AND_WO_3/w_0_0# gnd! 1.0fF
C75 m1_n188_6# gnd! 7.6fF
C76 PropagateGenerate_WO_0/2AND_WO_1/w_0_0# gnd! 1.0fF
C77 m2_189_369# gnd! 21.1fF
C78 PropagateGenerate_WO_0/XOR_WO_0/w_50_21# gnd! 2.7fF
C79 PropagateGenerate_WO_0/XOR_WO_0/a_51_n59# gnd! 1.6fF
C80 m2_n105_247# gnd! 4.6fF
C81 PropagateGenerate_WO_0/XOR_WO_1/w_50_21# gnd! 2.7fF
C82 PropagateGenerate_WO_0/XOR_WO_1/a_51_n59# gnd! 1.6fF
C83 m2_n89_397# gnd! 5.0fF
C84 m2_106_663# gnd! 24.4fF
C85 PropagateGenerate_WO_0/XOR_WO_2/w_50_21# gnd! 2.7fF
C86 PropagateGenerate_WO_0/XOR_WO_2/a_51_n59# gnd! 1.6fF
C87 m1_n193_459# gnd! 5.2fF
C88 m2_105_807# gnd! 25.9fF
C89 PropagateGenerate_WO_0/XOR_WO_3/w_50_21# gnd! 2.7fF
C90 PropagateGenerate_WO_0/XOR_WO_3/a_51_n59# gnd! 1.6fF
C91 m1_195_305# gnd! 2.1fF
C92 Carry_WO_0/w_7_77# gnd! 1.0fF
C93 Carry_WO_0/w_38_n91# gnd! 1.8fF
C94 Carry_WO_0/2NAND_WO_1/w_0_0# gnd! 1.0fF
C95 Carry_WO_0/m1_174_23# gnd! 1.2fF
C96 Carry_WO_0/3NAND_WO_0/w_0_0# gnd! 1.3fF
C97 m1_240_112# gnd! 14.9fF
C98 Carry_WO_0/2NAND_WO_2/w_0_0# gnd! 1.0fF
C99 Carry_WO_0/m1_395_n85# gnd! 1.5fF
C100 m1_240_299# gnd! 16.9fF
C101 Carry_WO_0/3NAND_WO_1/w_0_0# gnd! 1.3fF
C102 Carry_WO_0/m1_402_n83# gnd! 1.9fF
C103 Carry_WO_0/3NOR_WO_0/w_1_n3# gnd! 3.1fF
C104 m1_1395_46# gnd! 19.4fF
C105 m2_106_520# gnd! 26.6fF
C106 Carry_WO_0/4NAND_WO_0/w_0_0# gnd! 1.7fF
C107 Carry_WO_0/m1_409_n82# gnd! 4.6fF
C108 m1_243_38# gnd! 15.8fF
C109 Carry_WO_0/4NOR_WO_0/w_0_0# gnd! 4.6fF
C110 m1_1983_14# gnd! 5.9fF
C111 SUM_WO_0/XOR_WO_0/w_50_21# gnd! 2.7fF
C112 SUM_WO_0/XOR_WO_0/a_51_n59# gnd! 1.6fF
C113 m1_1978_186# gnd! 5.8fF
C114 SUM_WO_0/XOR_WO_1/w_50_21# gnd! 2.7fF
C115 SUM_WO_0/XOR_WO_1/a_51_n59# gnd! 1.6fF
C116 m1_1978_339# gnd! 5.6fF
C117 SUM_WO_0/XOR_WO_2/w_50_21# gnd! 2.7fF
C118 SUM_WO_0/XOR_WO_2/a_51_n59# gnd! 1.6fF
C119 m1_603_147# gnd! 7.5fF
C120 m1_1939_499# gnd! 5.3fF
C121 SUM_WO_0/XOR_WO_3/w_50_21# gnd! 2.7fF
C122 SUM_WO_0/XOR_WO_3/a_51_n59# gnd! 1.6fF
C123 m1_773_184# gnd! 7.3fF
C124 m1_1960_615# gnd! 2.4fF
C125 vdd gnd! 88.3fF
C126 m1_1015_205# gnd! 7.3fF
C127 FlipFlop_WO_0/w_0_0# gnd! 9.4fF
C128 FlipFlop_WO_1/w_0_0# gnd! 9.4fF
C129 FlipFlop_WO_2/w_0_0# gnd! 9.4fF
C130 FlipFlop_WO_3/w_0_0# gnd! 9.4fF
C131 a1 gnd! 3.8fF
C132 FlipFlop_WO_11/w_0_0# gnd! 9.4fF
C133 FlipFlop_WO_12/w_0_0# gnd! 9.4fF
C134 FlipFlop_WO_4/w_0_0# gnd! 9.4fF
