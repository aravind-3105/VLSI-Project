* SPICE3 file created from FlipFlop_WI.ext - technology: scmos

.option scale=0.09u

M1000 J1 D vdd w_0_0# pfet w=40 l=2
+  ad=240 pd=92 as=840 ps=362
M1001 J2 clk J1 w_0_0# pfet w=40 l=2
+  ad=560 pd=108 as=0 ps=0
M1002 J3 clk vdd w_0_0# pfet w=40 l=2
+  ad=680 pd=114 as=0 ps=0
M1003 Q_bar J3 vdd w_0_0# pfet w=40 l=2
+  ad=840 pd=202 as=0 ps=0
M1004 Q_bar vdd vdd w_0_0# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 Q Q_bar a_143_6# w_0_0# pfet w=40 l=2
+  ad=280 pd=94 as=280 ps=94
M1006 J2 D gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=500 ps=210
M1007 J4 clk gnd Gnd nfet w=20 l=2
+  ad=160 pd=56 as=0 ps=0
M1008 J3 J2 J4 Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1009 J5 J3 gnd Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1010 Q_bar a_94_n27# J5 Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1011 Q Q_bar gnd Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
C0 vdd w_0_0# 1.3fF
C1 clk gnd! 1.1fF
C2 w_0_0# gnd! 9.4fF
