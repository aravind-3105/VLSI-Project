magic
tech scmos
timestamp 1619596156
<< metal1 >>
rect 33 80 42 83
rect 39 72 42 80
rect 39 67 47 72
rect 1 37 9 41
rect 1 30 18 34
rect 28 30 51 34
rect 58 24 68 28
rect 27 0 68 3
use 2NAND_WO  2NAND_WO_0
timestamp 1619444932
transform 1 0 1 0 1 50
box -1 -50 32 33
use 2INV  2INV_0
timestamp 1619542334
transform 1 0 44 0 1 -44
box 0 45 24 116
<< labels >>
rlabel metal1 3 39 3 39 3 A
rlabel metal1 3 32 3 32 3 B
rlabel metal1 41 32 41 32 1 out_bar
rlabel metal1 66 26 66 26 7 out
rlabel metal1 38 1 38 1 1 gnd
rlabel metal1 41 82 41 82 5 vdd
<< end >>
