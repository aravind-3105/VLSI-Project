* SPICE3 file created from XOR.ext - technology: scmos

.option scale=0.09u

M1000 a_bar A vdd w_n1_0# pfet w=20 l=2
+  ad=100 pd=50 as=400 ps=200
M1001 a_30_6# a_bar vdd w_n1_0# pfet w=20 l=2
+  ad=160 pd=56 as=0 ps=0
M1002 out B a_30_6# w_n1_0# pfet w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M1003 a_66_6# a_43_n12# out w_n1_0# pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1004 vdd b_bar a_66_6# w_n1_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 vdd B b_bar w_n1_0# pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1006 a_bar A gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=200 ps=120
M1007 a_29_n32# B gnd Gnd nfet w=10 l=2
+  ad=160 pd=52 as=0 ps=0
M1008 out a_43_n12# a_29_n32# Gnd nfet w=10 l=2
+  ad=130 pd=66 as=0 ps=0
M1009 a_66_n32# a_bar out Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1010 gnd b_bar a_66_n32# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 gnd B b_bar Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50 ps=30
C0 a_bar gnd! 1.1fF
C1 w_n1_0# gnd! 4.5fF
