magic
tech scmos
timestamp 1619572441
<< metal1 >>
rect 58 172 358 176
rect 58 165 62 172
rect 206 165 210 172
rect 354 165 358 172
rect 154 121 156 125
rect 303 121 314 125
rect 145 29 154 33
rect 294 29 318 33
rect 0 0 412 4
<< m2contact >>
rect 149 121 154 126
rect 298 121 303 126
rect 121 78 126 83
rect 273 78 278 83
rect 420 78 425 83
rect 140 29 145 34
rect 289 29 294 34
<< metal2 >>
rect 121 -16 126 78
rect 140 34 145 189
rect 149 126 154 189
rect 273 -16 278 78
rect 289 34 294 189
rect 298 126 303 189
rect 420 -16 425 78
<< m345contact >>
rect 110 -22 427 -16
use XOR_WO  XOR_WO_0
timestamp 1619560144
transform 1 0 20 0 1 92
box -20 -92 103 77
use XOR_WO  XOR_WO_1
timestamp 1619560144
transform 1 0 172 0 1 92
box -20 -92 103 77
use XOR_WO  XOR_WO_2
timestamp 1619560144
transform 1 0 320 0 1 92
box -20 -92 103 77
<< end >>
