magic
tech scmos
timestamp 1619653108
<< metal1 >>
rect 21 701 26 731
rect 87 707 92 734
rect 113 701 118 731
rect 179 713 184 743
rect 325 604 526 609
rect 21 556 26 586
rect 87 562 92 589
rect 113 556 118 586
rect 179 563 184 593
rect 21 411 26 441
rect 87 417 92 444
rect 113 411 118 441
rect 179 420 184 450
rect 205 342 237 347
rect 195 305 212 309
rect 240 299 289 303
rect 21 265 26 295
rect 113 265 118 295
rect 205 259 237 264
rect 201 222 209 226
rect 325 220 329 604
rect 242 219 329 220
rect 219 216 329 219
rect 319 212 329 216
rect 205 155 237 160
rect 359 157 363 561
rect 294 153 363 157
rect 199 103 202 122
rect 240 112 319 116
rect 315 111 319 112
rect 409 111 413 561
rect 315 106 413 111
rect 167 81 237 86
rect 447 54 452 563
rect 1473 421 1560 426
rect 603 152 609 230
rect 773 189 778 215
rect 1015 210 1019 231
rect 1473 210 1478 421
rect 1015 205 1478 210
rect 1522 189 1527 354
rect 773 184 1527 189
rect 603 147 1553 152
rect 243 50 452 54
rect 1395 51 1400 112
rect 195 44 208 48
rect 243 38 246 50
rect 307 20 523 23
rect 224 18 523 20
rect 224 15 311 18
rect 1759 -14 1764 71
<< m2contact >>
rect 526 604 531 609
rect 289 298 294 303
rect 359 561 364 566
rect 409 561 414 566
rect 447 563 452 568
rect 289 153 294 158
rect 1560 421 1565 426
rect 1522 354 1527 359
rect 1553 147 1558 152
rect 1587 137 1592 142
rect 1395 112 1400 117
rect 1395 46 1400 51
rect 523 18 528 23
rect 1759 -19 1764 -14
<< metal2 >>
rect 301 811 530 814
rect 105 809 530 811
rect 105 807 307 809
rect 185 806 307 807
rect -124 687 -85 692
rect -124 678 -85 683
rect 307 667 474 670
rect 106 665 474 667
rect 106 663 310 665
rect 194 662 310 663
rect 470 638 474 665
rect 526 668 530 809
rect 526 663 625 668
rect 1362 663 1554 668
rect 516 653 529 658
rect 493 643 528 648
rect 470 633 723 638
rect 1366 633 1524 638
rect 364 623 590 628
rect 322 613 538 618
rect 1346 613 1500 618
rect -124 542 -85 547
rect -124 533 -85 538
rect 322 527 326 613
rect 1370 604 1395 609
rect 359 566 364 573
rect 409 566 414 573
rect 504 568 509 572
rect 452 564 509 568
rect 189 523 326 527
rect 106 522 326 523
rect 486 535 609 540
rect 106 520 311 522
rect 189 519 311 520
rect -124 397 -85 402
rect -124 384 -85 389
rect 189 372 425 377
rect 189 369 319 372
rect -124 247 -85 252
rect -124 231 -85 236
rect 289 158 294 298
rect 420 129 425 372
rect 486 142 490 535
rect 167 -32 172 4
rect 167 -33 173 -32
rect 486 -33 490 137
rect 524 23 528 467
rect 1496 219 1500 613
rect 1520 368 1524 633
rect 1548 515 1554 663
rect 1686 634 1780 639
rect 1548 510 1615 515
rect 1560 500 1625 505
rect 1560 426 1565 500
rect 1686 485 1780 490
rect 1520 363 1643 368
rect 1527 354 1579 359
rect 1686 338 1780 343
rect 1496 214 1643 219
rect 1553 205 1577 210
rect 1553 152 1558 205
rect 1686 186 1780 191
rect 563 137 1587 142
rect 538 60 543 124
rect 1395 117 1400 122
rect 538 55 1638 60
rect 1400 46 1735 51
rect 167 -53 490 -33
rect 524 -14 528 18
rect 582 -19 1759 -14
rect 524 -55 528 -19
<< m3contact >>
rect 511 653 516 658
rect 488 643 493 648
rect 359 623 364 628
rect 1395 604 1400 609
rect 359 573 364 578
rect 409 573 414 578
rect 504 572 509 577
rect 420 124 425 129
rect 486 137 491 142
rect 558 137 563 142
rect 538 124 543 129
rect 1395 122 1400 127
rect 524 -19 529 -14
rect 577 -19 582 -14
<< metal3 >>
rect 504 653 511 658
rect 409 643 488 648
rect 359 578 364 623
rect 409 578 414 643
rect 504 577 509 653
rect 491 137 558 142
rect 425 124 538 129
rect 1395 127 1400 604
rect 529 -19 577 -14
use PropagateGenerate_WO  PropagateGenerate_WO_0
timestamp 1619651442
transform 0 -1 184 1 0 251
box -254 -59 560 308
use Carry_WO  Carry_WO_0
timestamp 1619609411
transform 1 0 612 0 1 455
box -86 -250 759 213
use SUM_WO  SUM_WO_0
timestamp 1619592134
transform 0 -1 1764 1 0 65
box -19 -16 579 189
<< labels >>
rlabel metal2 417 -43 417 -43 1 vdd
rlabel metal2 526 -47 526 -47 1 gnd
rlabel metal1 606 207 606 207 1 c2
rlabel metal1 774 207 774 207 1 c3
rlabel metal1 1017 216 1017 216 1 c4
rlabel metal2 1773 188 1773 188 1 s1
rlabel metal2 1773 487 1773 487 1 s3
rlabel metal2 1771 637 1771 637 1 s4
rlabel metal2 1773 341 1773 341 1 s2
rlabel metal2 314 667 314 667 1 p3
rlabel metal1 323 51 323 51 1 g4
rlabel metal1 323 109 323 109 1 g3
rlabel metal1 320 155 320 155 1 g2
rlabel metal1 322 214 322 214 1 g1
rlabel metal2 314 524 314 524 1 p2
rlabel metal2 318 812 318 812 5 p4
rlabel metal1 200 111 200 111 1 g3_bar
rlabel metal1 202 47 202 47 1 g4_bar
rlabel metal1 204 224 204 224 1 g1_bar
rlabel metal1 200 307 200 307 1 g2_bar
rlabel metal2 -124 247 -85 252 1 a1
rlabel metal2 -124 231 -85 236 1 b1
rlabel metal2 -124 397 -85 402 1 a2
rlabel metal2 -124 542 -85 547 1 a3
rlabel metal2 -124 533 -85 538 1 b3
rlabel metal2 -124 687 -85 692 1 a4
rlabel metal2 -124 678 -85 683 1 b4
rlabel metal2 -124 384 -85 389 1 b2
<< end >>
