magic
tech scmos
timestamp 1619525138
<< metal1 >>
rect -121 204 172 210
rect -121 190 -115 204
rect 17 190 23 204
rect 166 192 172 204
rect -93 30 -21 35
rect 71 31 136 37
<< m2contact >>
rect -80 126 -73 133
rect 79 126 86 133
rect 237 128 244 135
rect -198 116 -191 122
rect -42 120 -35 126
rect 120 117 126 123
rect -199 76 -192 83
rect -41 79 -34 85
rect 117 80 124 86
<< metal2 >>
rect -243 2 -236 244
rect -225 83 -218 243
rect -206 122 -199 243
rect -206 116 -198 122
rect -225 76 -199 83
rect -78 2 -73 126
rect -62 85 -56 247
rect -47 126 -41 247
rect -47 120 -42 126
rect -62 79 -41 85
rect 80 3 86 126
rect 98 86 104 246
rect 113 123 119 246
rect 113 118 120 123
rect 114 117 120 118
rect 98 80 117 86
rect 238 5 244 128
use xor  xor_0
timestamp 1619522997
transform 1 0 -174 0 1 116
box -21 -87 98 78
use xor  xor_1
timestamp 1619522997
transform 1 0 -16 0 1 116
box -21 -87 98 78
use xor  xor_2
timestamp 1619522997
transform 1 0 143 0 1 118
box -21 -87 98 78
<< labels >>
rlabel metal2 -240 239 -240 239 3 p1
rlabel metal2 -240 13 -240 13 3 s1
rlabel metal2 -75 12 -75 12 1 s2
rlabel metal2 83 15 83 15 1 s3
rlabel metal2 241 17 241 17 7 s4
rlabel metal2 116 237 116 237 1 c3
rlabel metal2 101 236 101 236 1 p4
rlabel metal2 -44 239 -44 239 1 c2
rlabel metal2 -59 239 -59 239 1 p3
rlabel metal2 -222 237 -222 237 1 p2
rlabel metal2 -203 237 -203 237 1 c1
rlabel metal1 -59 32 -59 32 1 gnd
rlabel metal1 21 208 21 208 1 vdd
<< end >>
