.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.param W = {10*LAMBDA}
.param width_N={10*LAMBDA}
.param width_P={20*LAMBDA}
.global gnd vdd

Vdd	vdd	gnd	'SUPPLY'
vdA1     a1_d     0 pulse 0 0 0ns 100ps 100ps 5ns  30ns
vdA2     a2_d     0 pulse 1.8 0 0ns 100ps 100ps 30ns  30ns
vdA3     a3_d     0 pulse 0 0 0ns 100ps 100ps 10ns  30ns
vdA4     a4_d     0 pulse 1.8 0 0ns 100ps 100ps 30ns  30ns

vdB1     b1_d     0 pulse 0 0 0ns 100ps 100ps 10ns  30ns
vdB2     b2_d     0 pulse 0 0 0ns 100ps 100ps 10ns  30ns
vdB3     b3_d     0 pulse 1.8 0 0ns 100ps 100ps 30ns  30ns

vdB4     b4_d     0 pulse 1.8 0 0ns 100ps 100ps 30ns  30ns
* vdA1     a1_d     gnd 0   
* vdA2     a2_d     gnd 1.8
* vdA3     a3_d     gnd 0   
* vdA4     a4_d     gnd 1.8 

* vdB1     b1_d     gnd 0   
* vdB2     b2_d     gnd 0  
* vdB3     b3_d     gnd 1.8 
* vdB4     b4_d     gnd 1.8

vdC Ci 0 pulse 0 0 0ns 100ps 100ps 20ns 60ns
vclk   clk   0 pulse 0   1.8 0ns 100ps 100ps 20ns  40ns

.subckt xor_subckt a b y vdd gnd
//Top inverter
M1      a_bar       a       vdd     vdd  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
M2      a_bar       a       gnd     gnd  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

//Bottom Inverter
M3      b_bar       b       vdd     vdd  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
M4      b_bar       b       gnd     gnd  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

//Layer 2
M5      J1   a_bar    vdd     vdd  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
M6      y       b       J1     J1  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
M7      y       a       J2     J2  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
M8      J2      b     gnd     gnd  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

//Layer 3
M9      J11       b_bar    vdd     vdd  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
M10      y       a         J11     J11  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
M11      y     a_bar       J22     J22  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
M12      J22     b_bar     gnd     gnd  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
.ends xor_subckt


.subckt and_subckt a b y vdd gnd
.param w_AND_P = {2*W}
.param w_AND_N = {2*W}
* Layer-1
M1      nand       b       vdd     vdd  CMOSP   W={w_AND_P}   L={2*LAMBDA}
+ AS={5*w_AND_P*LAMBDA} PS={10*LAMBDA+2*w_AND_P} AD={5*w_AND_P*LAMBDA} PD={10*LAMBDA+2*w_AND_P}
M2      nand       a       vdd     vdd  CMOSP   W={w_AND_P}   L={2*LAMBDA}
+ AS={5*w_AND_P*LAMBDA} PS={10*LAMBDA+2*w_AND_P} AD={5*w_AND_P*LAMBDA} PD={10*LAMBDA+2*w_AND_P}
M3      nand       a       J     J  CMOSN   W={w_AND_N}   L={2*LAMBDA}
+ AS={5*w_AND_N*LAMBDA} PS={10*LAMBDA+2*w_AND_N} AD={5*w_AND_N*LAMBDA} PD={10*LAMBDA+2*w_AND_N}
M4      J         b      gnd gnd   CMOSN   W={w_AND_N}   L={2*LAMBDA}
+ AS={5*w_AND_N*LAMBDA} PS={10*LAMBDA+2*w_AND_N} AD={5*w_AND_N*LAMBDA} PD={10*LAMBDA+2*w_AND_N}

M5      y       nand       vdd     vdd  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
M6      y       nand       gnd     gnd  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
.ends and_subckt

.subckt or_subckt a b y vdd gnd
.param w_OR_P = {4*W}
.param w_OR_N = {W}
* Layer-1
M1      J1       a       vdd     vdd  CMOSP   W={w_OR_P}   L={2*LAMBDA}
+ AS={5*w_OR_P*LAMBDA} PS={10*LAMBDA+2*w_OR_P} AD={5*w_OR_P*LAMBDA} PD={10*LAMBDA+2*w_OR_P}
M2      nor      b       J1      J1  CMOSP   W={w_OR_P}   L={2*LAMBDA}
+ AS={5*w_OR_P*LAMBDA} PS={10*LAMBDA+2*w_OR_P} AD={5*w_OR_P*LAMBDA} PD={10*LAMBDA+2*w_OR_P}
M3      nor       a     gnd   gnd   CMOSN   W={w_OR_N}   L={2*LAMBDA}
+ AS={5*w_OR_N*LAMBDA} PS={10*LAMBDA+2*w_OR_N} AD={5*w_OR_N*LAMBDA} PD={10*LAMBDA+2*w_OR_N}
M4      nor       b     gnd   gnd   CMOSN   W={w_OR_N}   L={2*LAMBDA}
+ AS={5*w_OR_N*LAMBDA} PS={10*LAMBDA+2*w_OR_N} AD={5*w_OR_N*LAMBDA} PD={10*LAMBDA+2*w_OR_N}

M5      y       nor       vdd     vdd  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
M6      y       nor       gnd     gnd  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
.ends or_subckt

.subckt or3_subckt a b c y vdd gnd
.param w_OR_P3 = {6*W}
.param w_OR_N3 = {W}
// NOR
M1      J1       a       vdd     vdd  CMOSP   W={w_OR_P3}   L={2*LAMBDA}
+ AS={5*w_OR_P3*LAMBDA} PS={10*LAMBDA+2*w_OR_P3} AD={5*w_OR_P3*LAMBDA} PD={10*LAMBDA+2*w_OR_P3}

M2      J2       b       J1      J1  CMOSP   W={w_OR_P3}   L={2*LAMBDA}
+ AS={5*w_OR_P3*LAMBDA} PS={10*LAMBDA+2*w_OR_P3} AD={5*w_OR_P3*LAMBDA} PD={10*LAMBDA+2*w_OR_P3}

M3      nor      c       J2      J2  CMOSP   W={w_OR_P3}   L={2*LAMBDA}
+ AS={5*w_OR_P3*LAMBDA} PS={10*LAMBDA+2*w_OR_P3} AD={5*w_OR_P3*LAMBDA} PD={10*LAMBDA+2*w_OR_P3}

M4      nor       a     gnd   gnd   CMOSN   W={w_OR_N3}   L={2*LAMBDA}
+ AS={5*w_OR_N3*LAMBDA} PS={10*LAMBDA+2*w_OR_N3} AD={5*w_OR_N3*LAMBDA} PD={10*LAMBDA+2*w_OR_N3}

M5      nor       b     gnd   gnd   CMOSN   W={w_OR_N3}   L={2*LAMBDA}
+ AS={5*w_OR_N3*LAMBDA} PS={10*LAMBDA+2*w_OR_N3} AD={5*w_OR_N3*LAMBDA} PD={10*LAMBDA+2*w_OR_N3}

M6      nor       c     gnd   gnd   CMOSN   W={w_OR_N3}   L={2*LAMBDA}
+ AS={5*w_OR_N3*LAMBDA} PS={10*LAMBDA+2*w_OR_N3} AD={5*w_OR_N3*LAMBDA} PD={10*LAMBDA+2*w_OR_N3}

// Inverter
M7      y       nor       vdd     vdd  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

M8      y       nor       gnd     gnd  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
.ends or3_subckt

.subckt or4_subckt a b c d y vdd gnd
.param w_OR_P4 = {8*W}
.param w_OR_N4 = {W}
// NOR
M1      J1       a       vdd     vdd  CMOSP   W={w_OR_P4}   L={2*LAMBDA}
+ AS={5*w_OR_P4*LAMBDA} PS={10*LAMBDA+2*w_OR_P4} AD={5*w_OR_P4*LAMBDA} PD={10*LAMBDA+2*w_OR_P4}

M2      J2       b       J1      J1  CMOSP   W={w_OR_P4}   L={2*LAMBDA}
+ AS={5*w_OR_P4*LAMBDA} PS={10*LAMBDA+2*w_OR_P4} AD={5*w_OR_P4*LAMBDA} PD={10*LAMBDA+2*w_OR_P4}

M3      J3       c       J2      J2  CMOSP   W={w_OR_P4}   L={2*LAMBDA}
+ AS={5*w_OR_P4*LAMBDA} PS={10*LAMBDA+2*w_OR_P4} AD={5*w_OR_P4*LAMBDA} PD={10*LAMBDA+2*w_OR_P4}

M4      nor      d       J3      J3  CMOSP   W={w_OR_P4}   L={2*LAMBDA}
+ AS={5*w_OR_P4*LAMBDA} PS={10*LAMBDA+2*w_OR_P4} AD={5*w_OR_P4*LAMBDA} PD={10*LAMBDA+2*w_OR_P4}

M5      nor       a     gnd   gnd   CMOSN   W={w_OR_N4}   L={2*LAMBDA}
+ AS={5*w_OR_N4*LAMBDA} PS={10*LAMBDA+2*w_OR_N4} AD={5*w_OR_N4*LAMBDA} PD={10*LAMBDA+2*w_OR_N4}

M6      nor       b     gnd   gnd   CMOSN   W={w_OR_N4}   L={2*LAMBDA}
+ AS={5*w_OR_N4*LAMBDA} PS={10*LAMBDA+2*w_OR_N4} AD={5*w_OR_N4*LAMBDA} PD={10*LAMBDA+2*w_OR_N4}

M7      nor       c     gnd   gnd   CMOSN   W={w_OR_N4}   L={2*LAMBDA}
+ AS={5*w_OR_N4*LAMBDA} PS={10*LAMBDA+2*w_OR_N4} AD={5*w_OR_N4*LAMBDA} PD={10*LAMBDA+2*w_OR_N4}

M8      nor       d     gnd   gnd   CMOSN   W={w_OR_N4}   L={2*LAMBDA}
+ AS={5*w_OR_N4*LAMBDA} PS={10*LAMBDA+2*w_OR_N4} AD={5*w_OR_N4*LAMBDA} PD={10*LAMBDA+2*w_OR_N4}

// Inverter
M9      y       nor       vdd     vdd  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

M10      y       nor       gnd     gnd  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
.ends or4_subckt

.subckt and3_subckt a b c y vdd gnd
.param w_AND_P3 = {2*W}
.param w_AND_N3 = {3*W}
//NAND
M1      nand       a       vdd    vdd  CMOSP   W={w_AND_P3}   L={2*LAMBDA}
+ AS={5*w_AND_P3*LAMBDA} PS={10*LAMBDA+2*w_AND_P3} AD={5*w_AND_P3*LAMBDA} PD={10*LAMBDA+2*w_AND_P3}

M2      nand       b       vdd    vdd  CMOSP   W={w_AND_P3}   L={2*LAMBDA}
+ AS={5*w_AND_P3*LAMBDA} PS={10*LAMBDA+2*w_AND_P3} AD={5*w_AND_P3*LAMBDA} PD={10*LAMBDA+2*w_AND_P3}

M3      nand       c       vdd    vdd  CMOSP   W={w_AND_P3}   L={2*LAMBDA}
+ AS={5*w_AND_P3*LAMBDA} PS={10*LAMBDA+2*w_AND_P3} AD={5*w_AND_P3*LAMBDA} PD={10*LAMBDA+2*w_AND_P3}

M4      nand       a       J1     J1   CMOSN   W={w_AND_N3}   L={2*LAMBDA}
+ AS={5*w_AND_N3*LAMBDA} PS={10*LAMBDA+2*w_AND_N3} AD={5*w_AND_N3*LAMBDA} PD={10*LAMBDA+2*w_AND_N3}

M5      J1         b       J2     J2   CMOSN   W={w_AND_N3}   L={2*LAMBDA}
+ AS={5*w_AND_N3*LAMBDA} PS={10*LAMBDA+2*w_AND_N3} AD={5*w_AND_N3*LAMBDA} PD={10*LAMBDA+2*w_AND_N3}

M6      J2         c      gnd    gnd   CMOSN   W={w_AND_N3}   L={2*LAMBDA}
+ AS={5*w_AND_N3*LAMBDA} PS={10*LAMBDA+2*w_AND_N3} AD={5*w_AND_N3*LAMBDA} PD={10*LAMBDA+2*w_AND_N3}

//Inverter
M7      y       nand       vdd     vdd  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

M8      y       nand       gnd     gnd  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
.ends and3_subckt

.subckt and4_subckt a b c d y vdd gnd
.param w_AND_P4 = {2*W}
.param w_AND_N4 = {4*W}
//NAND
M1      nand       a       vdd    vdd  CMOSP   W={w_AND_P4}   L={2*LAMBDA}
+ AS={5*w_AND_P4*LAMBDA} PS={10*LAMBDA+2*w_AND_P4} AD={5*w_AND_P4*LAMBDA} PD={10*LAMBDA+2*w_AND_P4}

M2      nand       b       vdd    vdd  CMOSP   W={w_AND_P4}   L={2*LAMBDA}
+ AS={5*w_AND_P4*LAMBDA} PS={10*LAMBDA+2*w_AND_P4} AD={5*w_AND_P4*LAMBDA} PD={10*LAMBDA+2*w_AND_P4}

M3      nand       c       vdd    vdd  CMOSP   W={w_AND_P4}   L={2*LAMBDA}
+ AS={5*w_AND_P4*LAMBDA} PS={10*LAMBDA+2*w_AND_P4} AD={5*w_AND_P4*LAMBDA} PD={10*LAMBDA+2*w_AND_P4}

M4      nand       d       vdd    vdd  CMOSP   W={w_AND_P4}   L={2*LAMBDA}
+ AS={5*w_AND_P4*LAMBDA} PS={10*LAMBDA+2*w_AND_P4} AD={5*w_AND_P4*LAMBDA} PD={10*LAMBDA+2*width_P}

M5      nand       a       J1     J1   CMOSN   W={w_AND_N4}   L={2*LAMBDA}
+ AS={5*w_AND_N4*LAMBDA} PS={10*LAMBDA+2*w_AND_N4} AD={5*w_AND_N4*LAMBDA} PD={10*LAMBDA+2*w_AND_N4}

M6      J1         b       J2     J2   CMOSN   W={w_AND_N4}   L={2*LAMBDA}
+ AS={5*w_AND_N4*LAMBDA} PS={10*LAMBDA+2*w_AND_N4} AD={5*w_AND_N4*LAMBDA} PD={10*LAMBDA+2*w_AND_N4}

M7      J2         c       J3     J3   CMOSN   W={w_AND_N4}   L={2*LAMBDA}
+ AS={5*w_AND_N4*LAMBDA} PS={10*LAMBDA+2*w_AND_N4} AD={5*w_AND_N4*LAMBDA} PD={10*LAMBDA+2*w_AND_N4}

M8      J3         d      gnd    gnd   CMOSN   W={w_AND_N4}   L={2*LAMBDA}
+ AS={5*w_AND_N4*LAMBDA} PS={10*LAMBDA+2*w_AND_N4} AD={5*w_AND_N4*LAMBDA} PD={10*LAMBDA+2*w_AND_N4}

//Inverter
M9      y       nand       vdd     vdd  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

M10     y       nand       gnd     gnd  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
.ends and4_subckt


.subckt FlipFlop d clk q vdd gnd
// Layer-1
M1      J1       d       vdd     vdd  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

M2      J2       clk       J1     J1  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

M3      J2       d       gnd     gnd  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
// Layer-2
M4      J3       clk     vdd     vdd  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

M5      J3       J2        J4     J4  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

M6      J4       clk     gnd     gnd  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
// Layer-3
M7      q_bar     J3     vdd     vdd  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

M8      q_bar     clk      J5     J5  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

M9      J5        J3     gnd     gnd  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
// Layer-4
M10     q_bar     vdd    vdd     vdd  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
// Layer-5
M11      q       q_bar   vdd     vdd  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
M12      q       q_bar   gnd     gnd  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
.ends FlipFlop

xy11 a1_d clk a1 vdd gnd FlipFlop
xy21 a2_d clk a2 vdd gnd FlipFlop
xy12 a3_d clk a3 vdd gnd FlipFlop
xy22 a4_d clk a4 vdd gnd FlipFlop

xy13 b1_d clk b1 vdd gnd FlipFlop
xy23 b2_d clk b2 vdd gnd FlipFlop
xy14 b3_d clk b3 vdd gnd FlipFlop
xy24 b4_d clk b4 vdd gnd FlipFlop

// Propagate 
x1 a1 b1 P1 vdd gnd xor_subckt
x2 a2 b2 P2 vdd gnd xor_subckt
x3 a3 b3 P3 vdd gnd xor_subckt
x4 a4 b4 P4 vdd gnd xor_subckt

// Generate
x5 a1 b1 G1 vdd gnd and_subckt
x6 a2 b2 G2 vdd gnd and_subckt
x7 a3 b3 G3 vdd gnd and_subckt
x8 a4 b4 G4 vdd gnd and_subckt

// Carry Calculation
    // Cout1
    // Cout2
        x9  P2 G1 T2_1 vdd gnd and_subckt
        x10 G2 T2_1 Cout2 vdd gnd or_subckt
    // Cout3
        x11 P3 G2 T3_1 vdd gnd and_subckt
        x12 P3 P2 G1 T3_2 vdd gnd and3_subckt
        x13 G3 T3_1 T3_2 Cout3 vdd gnd or3_subckt
    // Cout4
        x14 P4 G3 T4_1 vdd gnd and_subckt
        x15 P4 P3 G2 T4_2 vdd gnd and3_subckt
        x16 P4 P3 P2 G1 T4_3 vdd gnd and4_subckt
        x17 G4 T4_1 T4_2 T4_3 Cout4 vdd gnd or4_subckt

// Sum 
x18 P1  Ci   Sum1 vdd gnd xor_subckt
x19 P2  G1   Sum2 vdd gnd xor_subckt
x20 P3 Cout2 Sum3 vdd gnd xor_subckt
x21 P4 Cout3 Sum4 vdd gnd xor_subckt

xS1 Sum1 clk S1 vdd gnd FlipFlop
xS2 Sum2 clk S2 vdd gnd FlipFlop
xS3 Sum3 clk S3 vdd gnd FlipFlop
xS4 Sum4 clk S4 vdd gnd FlipFlop

xC4 Cout4 clk Co4 vdd gnd FlipFlop


.tran 1n 200n
.control
set hcopypscolor = 1
set color0=white
set color1=black

run
plot (v(a1)+(2*v(a2))+(4*v(a3))+(8*v(a4)))/1.8
plot (v(a1_d)+(2*v(a2_d))+(4*v(a3_d))+(8*v(a4_d)))/1.8
plot (v(b1)+(2*v(b2))+(4*v(b3))+(8*v(b4)))/1.8
plot (v(b1_d)+(2*v(b2_d))+(4*v(b3_d))+(8*v(b4_d)))/1.8
plot (v(Sum1)+(2*v(Sum2))+(4*v(Sum3))+(8*v(Sum4)))/1.8
plot (v(S1)+(2*v(S2))+(4*v(S3))+(8*v(S4)))/1.8
plot v(Cout4)/1.8
plot v(Co4)/1.8
plot v(clk)/1.8
set curplottitle= "Aravind Narayanan-2019102014"
.endc