magic
tech scmos
timestamp 1619591882
<< metal1 >>
rect 58 172 506 176
rect 58 165 62 172
rect 206 165 210 172
rect 354 165 358 172
rect 502 165 506 172
rect -5 121 3 125
rect 154 121 156 125
rect 303 121 314 125
rect 450 121 462 125
rect 559 79 569 83
rect -14 29 0 33
rect 145 29 154 33
rect 294 29 318 33
rect 440 29 467 33
rect 0 0 579 4
<< m2contact >>
rect -10 121 -5 126
rect 149 121 154 126
rect 298 121 303 126
rect 445 121 450 126
rect 121 78 126 83
rect 273 78 278 83
rect 420 78 425 83
rect 569 78 574 83
rect -19 29 -14 34
rect 140 29 145 34
rect 289 29 294 34
rect 435 29 440 34
<< metal2 >>
rect -19 34 -14 189
rect -10 126 -5 189
rect 121 -16 126 78
rect 140 34 145 189
rect 149 126 154 189
rect 273 -16 278 78
rect 289 34 294 189
rect 298 126 303 189
rect 420 -16 425 78
rect 435 34 440 189
rect 445 126 450 189
rect 569 -16 574 78
use XOR_WO  XOR_WO_0
timestamp 1619560144
transform 1 0 20 0 1 92
box -20 -92 103 77
use XOR_WO  XOR_WO_1
timestamp 1619560144
transform 1 0 172 0 1 92
box -20 -92 103 77
use XOR_WO  XOR_WO_2
timestamp 1619560144
transform 1 0 320 0 1 92
box -20 -92 103 77
use XOR_WO  XOR_WO_3
timestamp 1619560144
transform 1 0 468 0 1 92
box -20 -92 103 77
<< labels >>
rlabel metal2 124 -11 124 -11 1 sum0
rlabel metal2 275 -11 275 -11 1 sum1
rlabel metal2 -8 184 -8 184 5 i0
rlabel metal2 -16 184 -16 184 4 j0
rlabel metal2 152 185 152 185 5 i1
rlabel metal2 142 185 142 185 5 j1
rlabel metal2 438 183 438 183 1 j3
rlabel metal2 448 183 448 183 1 i3
rlabel metal2 292 185 292 185 5 j2
rlabel metal2 301 185 301 185 5 i2
rlabel metal2 571 -9 571 -9 1 sum3
rlabel metal2 423 -9 423 -9 1 sum2
rlabel metal1 283 174 283 174 1 vdd
rlabel metal1 287 2 287 2 1 gnd
<< end >>
