magic
tech scmos
timestamp 1619552151
<< nwell >>
rect 50 21 98 77
<< ntransistor >>
rect 61 -51 63 -41
rect 69 -51 71 -41
rect 77 -51 79 -41
rect 85 -51 87 -41
<< ptransistor >>
rect 61 27 63 67
rect 69 27 71 67
rect 77 27 79 67
rect 85 27 87 67
<< ndiffusion >>
rect 60 -51 61 -41
rect 63 -51 69 -41
rect 71 -51 72 -41
rect 76 -51 77 -41
rect 79 -51 85 -41
rect 87 -51 88 -41
<< pdiffusion >>
rect 60 27 61 67
rect 63 27 64 67
rect 68 27 69 67
rect 71 27 72 67
rect 76 27 77 67
rect 79 27 80 67
rect 84 27 85 67
rect 87 27 88 67
<< ndcontact >>
rect 56 -51 60 -41
rect 72 -51 76 -41
rect 88 -51 92 -41
<< pdcontact >>
rect 6 42 10 62
rect 56 27 60 67
rect 64 27 68 67
rect 72 27 76 67
rect 80 27 84 67
rect 88 27 92 67
<< polysilicon >>
rect 61 67 63 70
rect 69 67 71 70
rect 77 67 79 70
rect 85 67 87 70
rect 61 -41 63 27
rect 69 11 71 27
rect 69 -41 71 7
rect 77 3 79 27
rect 77 -41 79 -1
rect 85 -26 87 27
rect 85 -41 87 -30
rect 61 -65 63 -51
rect 69 -65 71 -51
rect 77 -65 79 -51
rect 85 -65 87 -51
<< polycontact >>
rect 57 14 61 18
rect 67 7 71 11
rect 75 -1 79 3
rect 83 -30 87 -26
<< metal1 >>
rect 20 73 68 77
rect 20 71 24 73
rect -1 66 24 71
rect 64 67 68 73
rect -8 29 7 33
rect -8 -2 -4 29
rect 14 23 34 27
rect 72 73 92 77
rect 72 67 76 73
rect 88 67 92 73
rect 56 24 60 27
rect 72 24 76 27
rect 56 21 76 24
rect 43 14 57 18
rect 0 0 22 5
rect -15 -3 -4 -2
rect 43 -3 47 14
rect 80 11 84 27
rect -15 -7 47 -3
rect 50 7 67 11
rect 80 7 98 11
rect 50 -10 53 7
rect -15 -14 53 -10
rect 56 -1 75 3
rect -15 -59 -11 -14
rect 56 -18 60 -1
rect -1 -26 24 -21
rect 41 -30 83 -26
rect -15 -63 7 -59
rect 41 -65 45 -30
rect 90 -33 94 7
rect 72 -37 94 -33
rect 72 -41 76 -37
rect 14 -69 45 -65
rect 56 -87 60 -51
rect 88 -87 92 -51
rect -15 -92 24 -87
rect 29 -92 92 -87
<< m2contact >>
rect -6 66 -1 71
rect 34 23 39 28
rect 22 0 27 5
rect -6 -26 -1 -21
rect 55 -23 60 -18
rect 24 -92 29 -87
<< metal2 >>
rect -6 -21 -2 66
rect 23 -16 27 0
rect 23 -20 29 -16
rect 25 -87 29 -20
rect 35 -18 39 23
rect 35 -23 55 -18
use 2INV  2INV_0
timestamp 1619542334
transform 1 0 0 0 1 -45
box 0 45 24 116
use 2INV  2INV_1
timestamp 1619542334
transform 1 0 0 0 1 -137
box 0 45 24 116
<< labels >>
rlabel metal1 95 9 95 9 7 out
rlabel metal1 37 -91 37 -91 1 gnd
rlabel metal1 38 75 38 75 5 vdd
rlabel metal1 14 23 34 27 1 A_bar
rlabel metal1 0 -61 0 -61 1 B
rlabel metal1 19 -67 19 -67 1 B_bar
rlabel metal1 1 29 6 33 1 A
<< end >>
