magic
tech scmos
timestamp 1619595931
<< metal1 >>
rect 33 80 42 83
rect 39 72 42 80
rect 39 67 47 72
rect 29 30 49 34
rect 27 0 68 3
use 2NAND_WO  2NAND_WO_0
timestamp 1619444932
transform 1 0 1 0 1 50
box -1 -50 32 33
use 2INV  2INV_0
timestamp 1619542334
transform 1 0 44 0 1 -44
box 0 45 24 116
<< end >>
