* SPICE3 file created from GenProp_WI.ext - technology: scmos
.include TSMC_180nm.txt
.option scale=0.09u
.param SUPPLY=1.8
.param LAMBDA=0.09u
.global gnd vdd

Vdd	vdd	gnd	'SUPPLY'
vd1a a0  0 pulse 1.8 0 0ns 100ps 100ps 20ns  40ns
vd2a a1  0 pulse 1.8 0 0ns 100ps 100ps 50ns  80ns
vd3a a2  0 pulse 1.8 0 0ns 100ps 100ps 80ns  120ns
vd4a a3  0 pulse 1.8 0 0ns 100ps 100ps 160ns 320ns

vd1b b0  0 pulse 1.8 0 0ns 100ps 100ps 20ns  40ns
vd2b b1  0 pulse 1.8 0 0ns 100ps 100ps 40ns  80ns
vd3b b2  0 pulse 1.8 0 0ns 100ps 100ps 80ns  160ns
vd4b b3  0 pulse 1.8 0 0ns 100ps 100ps 160ns 320ns

M1000 XOR_WO_3/a_59_n30# b3 vdd XOR_WO_3/2INV_1/w_0_81# CMOSP w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1001 XOR_WO_3/a_59_n30# b3 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=1200 ps=680
M1002 XOR_WO_3/a_51_n59# a3 vdd XOR_WO_3/2INV_0/w_0_81# CMOSP w=20 l=2
+  ad=100 pd=50 as=2160 ps=968
M1003 XOR_WO_3/a_51_n59# a3 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1004 vdd XOR_WO_3/a_51_n59# XOR_WO_3/a_56_27# XOR_WO_3/w_50_21# CMOSP w=40 l=2
+  ad=0 pd=0 as=400 ps=180
M1005 XOR_WO_3/a_71_27# XOR_WO_3/a_59_n30# vdd XOR_WO_3/w_50_21# CMOSP w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1006 p3 a3 XOR_WO_3/a_71_27# XOR_WO_3/w_50_21# CMOSP w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1007 XOR_WO_3/a_56_27# b3 p3 XOR_WO_3/w_50_21# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1008 XOR_WO_3/a_63_n51# XOR_WO_3/a_59_n30# gnd gnd CMOSN w=10 l=2
+  ad=60 pd=32 as=0 ps=01.8 0
M1009 p3 XOR_WO_3/a_51_n59# XOR_WO_3/a_63_n51# gnd CMOSN w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1010 XOR_WO_3/a_79_n51# a3 p3 gnd CMOSN w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1011 gnd b3 XOR_WO_3/a_79_n51# gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1012 XOR_WO_2/a_59_n30# b2 vdd XOR_WO_2/2INV_1/w_0_81# CMOSP w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1013 XOR_WO_2/a_59_n30# b2 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1014 XOR_WO_2/a_51_n59# a2 vdd XOR_WO_2/2INV_0/w_0_81# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1015 XOR_WO_2/a_51_n59# a2 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1016 vdd XOR_WO_2/a_51_n59# XOR_WO_2/a_56_27# XOR_WO_2/w_50_21# CMOSP w=40 l=2
+  ad=0 pd=0 as=400 ps=180
M1017 XOR_WO_2/a_71_27# XOR_WO_2/a_59_n30# vdd XOR_WO_2/w_50_21# CMOSP w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1018 p2 a2 XOR_WO_2/a_71_27# XOR_WO_2/w_50_21# CMOSP w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1019 XOR_WO_2/a_56_27# b2 p2 XOR_WO_2/w_50_21# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1020 XOR_WO_2/a_63_n51# XOR_WO_2/a_59_n30# gnd gnd CMOSN w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1021 p2 XOR_WO_2/a_51_n59# XOR_WO_2/a_63_n51# gnd CMOSN w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1022 XOR_WO_2/a_79_n51# a2 p2 gnd CMOSN w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1023 gnd b2 XOR_WO_2/a_79_n51# gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1024 XOR_WO_1/a_59_n30# b1 vdd XOR_WO_1/2INV_1/w_0_81# CMOSP w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1025 XOR_WO_1/a_59_n30# b1 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1026 XOR_WO_1/a_51_n59# a1 vdd XOR_WO_1/2INV_0/w_0_81# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1027 XOR_WO_1/a_51_n59# a1 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1028 vdd XOR_WO_1/a_51_n59# XOR_WO_1/a_56_27# XOR_WO_1/w_50_21# CMOSP w=40 l=2
+  ad=0 pd=0 as=400 ps=180
M1029 XOR_WO_1/a_71_27# XOR_WO_1/a_59_n30# vdd XOR_WO_1/w_50_21# CMOSP w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1030 p1 a1 XOR_WO_1/a_71_27# XOR_WO_1/w_50_21# CMOSP w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1031 XOR_WO_1/a_56_27# b1 p1 XOR_WO_1/w_50_21# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1032 XOR_WO_1/a_63_n51# XOR_WO_1/a_59_n30# gnd gnd CMOSN w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1033 p1 XOR_WO_1/a_51_n59# XOR_WO_1/a_63_n51# gnd CMOSN w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1034 XOR_WO_1/a_79_n51# a1 p1 gnd CMOSN w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1035 gnd b1 XOR_WO_1/a_79_n51# gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0



M1036 XOR_WO_0/a_59_n30# b0 vdd XOR_WO_0/2INV_1/w_0_81# CMOSP w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1037 XOR_WO_0/a_59_n30# b0 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1038 XOR_WO_0/a_51_n59# a0 vdd XOR_WO_0/2INV_0/w_0_81# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1039 XOR_WO_0/a_51_n59# a0 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1040 vdd XOR_WO_0/a_51_n59# XOR_WO_0/a_56_27# XOR_WO_0/w_50_21# CMOSP w=40 l=2
+  ad=0 pd=0 as=400 ps=180
M1041 XOR_WO_0/a_71_27# XOR_WO_0/a_59_n30# vdd XOR_WO_0/w_50_21# CMOSP w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1042 p0 a0 XOR_WO_0/a_71_27# XOR_WO_0/w_50_21# CMOSP w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1043 XOR_WO_0/a_56_27# b0 p0 XOR_WO_0/w_50_21# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1044 XOR_WO_0/a_63_n51# XOR_WO_0/a_59_n30# gnd gnd CMOSN w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1045 p0 XOR_WO_0/a_51_n59# XOR_WO_0/a_63_n51# gnd CMOSN w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1046 XOR_WO_0/a_79_n51# a0 p0 gnd CMOSN w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1047 gnd b0 XOR_WO_0/a_79_n51# gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1048 g1_bar a1 vdd 2AND_WO_1/w_0_0# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1049 vdd b1 g1_bar 2AND_WO_1/w_0_0# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1050 2AND_WO_1/a_13_n43# a1 gnd gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1051 g1_bar b1 2AND_WO_1/a_13_n43# gnd CMOSN w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1052 g3_bar a3 vdd 2AND_WO_3/w_0_0# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1053 vdd b3 g3_bar 2AND_WO_3/w_0_0# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1054 2AND_WO_3/a_13_n43# a3 gnd gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1055 g3_bar b3 2AND_WO_3/a_13_n43# gnd CMOSN w=20 l=2
+  ad=140 pd=54 as=0 ps=0

M1056 g0_bar a0 vdd 2AND_WO_0/w_0_0# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1057 vdd b0 g0_bar 2AND_WO_0/w_0_0# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1058 2AND_WO_0/a_13_n43# a0 gnd gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1059 g0_bar b0 2AND_WO_0/a_13_n43# gnd CMOSN w=20 l=2
+  ad=140 pd=54 as=0 ps=0

M1060 g2_bar a2 vdd 2AND_WO_2/w_0_0# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1061 vdd b2 g2_bar 2AND_WO_2/w_0_0# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1062 2AND_WO_2/a_13_n43# a2 gnd gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1063 g2_bar b2 2AND_WO_2/a_13_n43# gnd CMOSN w=20 l=2
+  ad=140 pd=54 as=0 ps=0


M1064 g1 g1_bar vdd vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1065 g1 g1_bar gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=1400 ps=800
M1066 g0 g0_bar vdd 2INV_2/w_0_81# CMOSP w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1067 g0 g0_bar gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1068 g2 g2_bar vdd 2INV_1/w_0_81# CMOSP w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1069 g2 g2_bar gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1070 g3 g3_bar vdd 2INV_0/w_0_81# CMOSP w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1071 g3 g3_bar gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0


C0 XOR_WO_1/a_56_27# p1 1.1fF
C1 a0 b0 3.5fF
C2 a3 b2 5.2fF
C3 a1 b1 4.8fF
C4 a2 b2 7.4fF
C5 a3 b3 12.6fF
C6 vdd g0_bar 1.2fF
C7 XOR_WO_0/a_56_27# p0 1.1fF
C8 XOR_WO_2/a_56_27# p2 1.1fF
C9 XOR_WO_3/a_56_27# p3 1.1fF
C10 a2 b1 2.4fF
C11 g2_bar gnd 1.4fF
C12 b2 gnd 8.3fF
C13 2AND_WO_2/w_0_0# gnd 1.0fF
C14 gnd gnd 11.7fF
C15 g0_bar gnd 1.0fF
C16 b0 gnd 4.1fF
C17 2AND_WO_0/w_0_0# gnd 1.0fF
C18 b3 gnd 7.4fF
C19 2AND_WO_3/w_0_0# gnd 1.0fF
C20 b1 gnd 5.8fF
C21 2AND_WO_1/w_0_0# gnd 1.0fF
C22 p0 gnd 1.5fF
C23 XOR_WO_0/w_50_21# gnd 2.7fF
C24 XOR_WO_0/a_51_n59# gnd 1.6fF
C25 a0 gnd 3.5fF
C26 p1 gnd 1.5fF
C27 XOR_WO_1/w_50_21# gnd 2.7fF
C28 XOR_WO_1/a_51_n59# gnd 1.6fF
C29 a1 gnd 3.8fF
C30 p2 gnd 1.5fF
C31 XOR_WO_2/w_50_21# gnd 2.7fF
C32 XOR_WO_2/a_51_n59# gnd 1.6fF
C33 a2 gnd 6.9fF
C34 p3 gnd 1.5fF
C35 XOR_WO_3/w_50_21# gnd 2.7fF
C36 vdd gnd 1.7fF
C37 XOR_WO_3/a_51_n59# gnd 1.6fF
C38 a3 gnd 6.5fF
C39 g1_bar gnd 2.1fF


.tran 1n 320n
.control
set hcopypscolor = 1
set color0=white
set color1=black

run
set curplottitle= "Aravind Narayanan-2019102014"
plot v(a0)/1.8 ((v(b0)/1.8)+2) ((v(g0)/1.8)+4) ((v(p0)/1.8)+6)  
plot v(a1)/1.8 ((v(b1)/1.8)+2) ((v(g1)/1.8)+4) ((v(p1)/1.8)+6) 
plot v(a2)/1.8 ((v(b2)/1.8)+2) ((v(g2)/1.8)+4) ((v(p2)/1.8)+6) 
plot v(a3)/1.8 ((v(b3)/1.8)+2) ((v(g3)/1.8)+4) ((v(p3)/1.8)+6) 
.endc