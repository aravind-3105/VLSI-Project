magic
tech scmos
timestamp 1619640426
<< nwell >>
rect 0 53 148 57
rect 0 0 165 53
<< ntransistor >>
rect 11 -52 13 -32
rect 53 -52 55 -32
rect 63 -52 65 -32
rect 88 -52 90 -32
rect 96 -52 98 -32
rect 150 -52 152 -32
<< ptransistor >>
rect 11 6 13 46
rect 19 6 21 46
rect 53 6 55 46
rect 88 6 90 46
rect 123 6 125 46
rect 150 6 152 46
<< ndiffusion >>
rect 10 -52 11 -32
rect 13 -52 14 -32
rect 52 -52 53 -32
rect 55 -52 63 -32
rect 65 -52 68 -32
rect 84 -52 88 -32
rect 90 -52 96 -32
rect 98 -52 101 -32
rect 147 -52 150 -32
rect 152 -52 155 -32
<< pdiffusion >>
rect 10 6 11 46
rect 13 6 19 46
rect 21 6 31 46
rect 52 6 53 46
rect 55 6 68 46
rect 87 6 88 46
rect 90 6 101 46
rect 121 6 123 46
rect 125 6 127 46
rect 143 6 150 46
rect 152 6 155 46
<< ndcontact >>
rect 6 -52 10 -32
rect 14 -52 18 -32
rect 48 -52 52 -32
rect 68 -52 72 -32
rect 80 -52 84 -32
rect 101 -52 105 -32
rect 143 -52 147 -32
rect 155 -52 159 -32
<< pdcontact >>
rect 6 6 10 46
rect 31 6 35 46
rect 48 6 52 46
rect 68 6 72 46
rect 83 6 87 46
rect 101 6 105 46
rect 117 6 121 46
rect 127 6 131 46
rect 155 6 159 46
<< polysilicon >>
rect 11 46 13 49
rect 19 46 21 49
rect 53 46 55 50
rect 88 46 90 49
rect 123 46 125 49
rect 150 46 152 49
rect 11 -3 13 6
rect 11 -32 13 -7
rect 19 -10 21 6
rect 53 -2 55 6
rect 88 -4 90 6
rect 19 -18 21 -14
rect 53 -32 55 -6
rect 63 -32 65 -22
rect 88 -32 90 -8
rect 96 -32 98 -27
rect 123 -35 125 6
rect 150 -15 152 6
rect 150 -32 152 -19
rect 123 -41 125 -39
rect 11 -55 13 -52
rect 53 -55 55 -52
rect 63 -55 65 -52
rect 88 -55 90 -52
rect 96 -55 98 -52
rect 150 -57 152 -52
<< polycontact >>
rect 9 -7 13 -3
rect 51 -6 55 -2
rect 17 -14 21 -10
rect 86 -8 90 -4
rect 61 -22 65 -18
rect 94 -27 98 -23
rect 148 -19 152 -15
rect 121 -39 125 -35
<< metal1 >>
rect 0 53 109 57
rect 0 52 87 53
rect 114 53 165 57
rect 6 46 10 52
rect 48 46 52 52
rect 83 46 87 52
rect 117 46 121 53
rect 143 6 147 53
rect 0 -7 9 -3
rect -1 -14 17 -10
rect 21 -14 23 -10
rect 31 -18 35 6
rect 38 -6 51 -2
rect 68 -4 72 6
rect 38 -9 43 -6
rect 68 -8 86 -4
rect 31 -22 61 -18
rect 31 -28 35 -22
rect 14 -32 35 -28
rect 68 -32 72 -8
rect 76 -23 81 -17
rect 101 -15 105 6
rect 127 -15 131 6
rect 155 -5 159 6
rect 155 -9 165 -5
rect 101 -19 148 -15
rect 76 -27 94 -23
rect 101 -32 105 -19
rect 155 -32 159 -9
rect 116 -39 121 -35
rect 6 -59 10 -52
rect 48 -59 52 -52
rect 80 -59 84 -52
rect 143 -59 147 -52
rect 6 -64 164 -59
<< m2contact >>
rect 109 52 114 57
rect 23 -14 28 -9
rect 38 -14 43 -9
rect 76 -17 81 -12
rect 111 -39 116 -34
<< metal2 >>
rect 55 -6 65 -2
rect 28 -14 38 -10
rect 61 -12 65 -6
rect 61 -15 76 -12
rect 111 -34 114 52
<< labels >>
rlabel metal1 163 -7 163 -7 7 Q
rlabel metal1 110 -62 110 -62 1 gnd
rlabel metal1 99 55 99 55 5 vdd
rlabel metal1 3 -5 3 -5 3 D
rlabel metal1 3 -12 3 -12 3 clk
rlabel pdiffusion 16 25 16 25 1 J1
rlabel pdiffusion 26 25 26 25 1 J2
rlabel pdiffusion 60 27 60 27 1 J3
rlabel ndiffusion 59 -42 59 -42 1 J4
rlabel ndiffusion 93 -42 93 -42 1 J5
rlabel metal1 105 -16 105 -16 1 Q_bar
<< end >>
