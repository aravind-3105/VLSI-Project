.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.option scale=0.09u
.global gnd vdd



Vdd	vdd	gnd	'SUPPLY'
vd10     a1in     0 pulse 0 1.8 10ns 0ps 0ps 5ns  1600ns
vd_bar10 a1in_inv 0 pulse 1.8 0 10ns 0ps 0ps 5ns  1600ns

vd20    b1in     0 pulse 0 1.8 10ns 0ps 0ps 5ns  1600ns
vd_bar20 b1in_inv 0 pulse 1.8 0 10ns 0ps 0ps 5ns  1600ns

vd11     a2in     0 pulse 0 1.8 10ns 0ps 0ps 5ns  1600ns
vd_bar11 a2in_inv 0 pulse 1.8 0 10ns 0ps 0ps 5ns  1600ns

vd21     b2in     gnd 0
vd_bar21 b2in_inv vdd 0

vd12     a3in     0 pulse 0 1.8 10ns 0ps 0ps 5ns  1600ns
vd_bar12 a3in_inv 0 pulse 1.8 0 10ns 0ps 0ps 5ns  1600ns

vd22     b3in     gnd 0
vd_bar22 b3in_inv vdd 0

vd13     a4in     0 pulse 0 1.8 10ns 0ps 0ps 5ns  1600ns
vd_bar13 a4in_inv 0 pulse 1.8 0 10ns 0ps 0ps 5ns  1600ns

vd23     b4in     0 pulse 0 1.8 10ns 0ps 0ps 5ns  1600ns
vd_bar23 b4in_inv 0 pulse 1.8 0 10ns 0ps 0ps 5ns  1600ns

vclk   clk   0 pulse 0   1.8 0ns 0ps 0ps 20ns  40ns


M1000 s4out dff_12/dlatch_1/m1_29_n71# vdd dff_12/dlatch_1/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=30040 ps=14740
M1001 vdd m2_2425_n861# s4out dff_12/dlatch_1/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 dff_12/dlatch_1/nand_3/a_n33_20# dff_12/dlatch_1/m1_29_n71# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=14480 ps=7418
M1003 s4out m2_2425_n861# dff_12/dlatch_1/nand_3/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1004 dff_12/dlatch_1/m1_29_n71# clk vdd dff_12/dlatch_1/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1005 vdd dff_12/m1_n21_n58# dff_12/dlatch_1/m1_29_n71# dff_12/dlatch_1/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 dff_12/dlatch_1/nand_2/a_n33_20# clk gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1007 dff_12/dlatch_1/m1_29_n71# dff_12/m1_n21_n58# dff_12/dlatch_1/nand_2/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1008 m2_2425_n861# dff_12/dlatch_1/m1_27_49# vdd dff_12/dlatch_1/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1009 vdd s4out m2_2425_n861# dff_12/dlatch_1/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1010 dff_12/dlatch_1/nand_1/a_n33_20# dff_12/dlatch_1/m1_27_49# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1011 m2_2425_n861# s4out dff_12/dlatch_1/nand_1/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1012 dff_12/dlatch_1/m1_27_49# clk vdd dff_12/dlatch_1/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1013 vdd dff_12/m1_n9_n58# dff_12/dlatch_1/m1_27_49# dff_12/dlatch_1/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1014 dff_12/dlatch_1/nand_0/a_n33_20# clk gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1015 dff_12/dlatch_1/m1_27_49# dff_12/m1_n9_n58# dff_12/dlatch_1/nand_0/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1016 dff_12/m1_n21_n58# dff_12/dlatch_0/m1_29_n71# vdd dff_12/dlatch_0/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1017 vdd dff_12/m1_n9_n58# dff_12/m1_n21_n58# dff_12/dlatch_0/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1018 dff_12/dlatch_0/nand_3/a_n33_20# dff_12/dlatch_0/m1_29_n71# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1019 dff_12/m1_n21_n58# dff_12/m1_n9_n58# dff_12/dlatch_0/nand_3/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1020 dff_12/dlatch_0/m1_29_n71# dff_12/m1_n65_174# vdd dff_12/dlatch_0/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1021 vdd s4 dff_12/dlatch_0/m1_29_n71# dff_12/dlatch_0/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1022 dff_12/dlatch_0/nand_2/a_n33_20# dff_12/m1_n65_174# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1023 dff_12/dlatch_0/m1_29_n71# s4 dff_12/dlatch_0/nand_2/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1024 dff_12/m1_n9_n58# dff_12/dlatch_0/m1_27_49# vdd dff_12/dlatch_0/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1025 vdd dff_12/m1_n21_n58# dff_12/m1_n9_n58# dff_12/dlatch_0/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1026 dff_12/dlatch_0/nand_1/a_n33_20# dff_12/dlatch_0/m1_27_49# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1027 dff_12/m1_n9_n58# dff_12/m1_n21_n58# dff_12/dlatch_0/nand_1/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1028 dff_12/dlatch_0/m1_27_49# dff_12/m1_n65_174# vdd dff_12/dlatch_0/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1029 vdd s4_inv dff_12/dlatch_0/m1_27_49# dff_12/dlatch_0/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1030 dff_12/dlatch_0/nand_0/a_n33_20# dff_12/m1_n65_174# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1031 dff_12/dlatch_0/m1_27_49# s4_inv dff_12/dlatch_0/nand_0/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1032 dff_12/m1_n65_174# clk vdd dff_12/inv_0/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1033 dff_12/m1_n65_174# clk gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1034 s3out dff_11/dlatch_1/m1_29_n71# vdd dff_11/dlatch_1/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1035 vdd m2_1903_n872# s3out dff_11/dlatch_1/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1036 dff_11/dlatch_1/nand_3/a_n33_20# dff_11/dlatch_1/m1_29_n71# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1037 s3out m2_1903_n872# dff_11/dlatch_1/nand_3/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1038 dff_11/dlatch_1/m1_29_n71# clk vdd dff_11/dlatch_1/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1039 vdd dff_11/m1_n21_n58# dff_11/dlatch_1/m1_29_n71# dff_11/dlatch_1/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1040 dff_11/dlatch_1/nand_2/a_n33_20# clk gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1041 dff_11/dlatch_1/m1_29_n71# dff_11/m1_n21_n58# dff_11/dlatch_1/nand_2/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1042 m2_1903_n872# dff_11/dlatch_1/m1_27_49# vdd dff_11/dlatch_1/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1043 vdd s3out m2_1903_n872# dff_11/dlatch_1/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1044 dff_11/dlatch_1/nand_1/a_n33_20# dff_11/dlatch_1/m1_27_49# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1045 m2_1903_n872# s3out dff_11/dlatch_1/nand_1/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1046 dff_11/dlatch_1/m1_27_49# clk vdd dff_11/dlatch_1/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1047 vdd dff_11/m1_n9_n58# dff_11/dlatch_1/m1_27_49# dff_11/dlatch_1/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1048 dff_11/dlatch_1/nand_0/a_n33_20# clk gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1049 dff_11/dlatch_1/m1_27_49# dff_11/m1_n9_n58# dff_11/dlatch_1/nand_0/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1050 dff_11/m1_n21_n58# dff_11/dlatch_0/m1_29_n71# vdd dff_11/dlatch_0/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1051 vdd dff_11/m1_n9_n58# dff_11/m1_n21_n58# dff_11/dlatch_0/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1052 dff_11/dlatch_0/nand_3/a_n33_20# dff_11/dlatch_0/m1_29_n71# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1053 dff_11/m1_n21_n58# dff_11/m1_n9_n58# dff_11/dlatch_0/nand_3/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1054 dff_11/dlatch_0/m1_29_n71# dff_11/m1_n65_174# vdd dff_11/dlatch_0/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1055 vdd s3 dff_11/dlatch_0/m1_29_n71# dff_11/dlatch_0/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1056 dff_11/dlatch_0/nand_2/a_n33_20# dff_11/m1_n65_174# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1057 dff_11/dlatch_0/m1_29_n71# s3 dff_11/dlatch_0/nand_2/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1058 dff_11/m1_n9_n58# dff_11/dlatch_0/m1_27_49# vdd dff_11/dlatch_0/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1059 vdd dff_11/m1_n21_n58# dff_11/m1_n9_n58# dff_11/dlatch_0/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1060 dff_11/dlatch_0/nand_1/a_n33_20# dff_11/dlatch_0/m1_27_49# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1061 dff_11/m1_n9_n58# dff_11/m1_n21_n58# dff_11/dlatch_0/nand_1/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1062 dff_11/dlatch_0/m1_27_49# dff_11/m1_n65_174# vdd dff_11/dlatch_0/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1063 vdd m1_1732_n280# dff_11/dlatch_0/m1_27_49# dff_11/dlatch_0/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1064 dff_11/dlatch_0/nand_0/a_n33_20# dff_11/m1_n65_174# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1065 dff_11/dlatch_0/m1_27_49# m1_1732_n280# dff_11/dlatch_0/nand_0/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1066 dff_11/m1_n65_174# clk vdd dff_11/inv_0/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1067 dff_11/m1_n65_174# clk gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1068 s2out dff_10/dlatch_1/m1_29_n71# vdd dff_10/dlatch_1/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1069 vdd m2_1376_n866# s2out dff_10/dlatch_1/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1070 dff_10/dlatch_1/nand_3/a_n33_20# dff_10/dlatch_1/m1_29_n71# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1071 s2out m2_1376_n866# dff_10/dlatch_1/nand_3/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1072 dff_10/dlatch_1/m1_29_n71# clk vdd dff_10/dlatch_1/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1073 vdd dff_10/m1_n21_n58# dff_10/dlatch_1/m1_29_n71# dff_10/dlatch_1/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1074 dff_10/dlatch_1/nand_2/a_n33_20# clk gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1075 dff_10/dlatch_1/m1_29_n71# dff_10/m1_n21_n58# dff_10/dlatch_1/nand_2/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1076 m2_1376_n866# dff_10/dlatch_1/m1_27_49# vdd dff_10/dlatch_1/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1077 vdd s2out m2_1376_n866# dff_10/dlatch_1/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1078 dff_10/dlatch_1/nand_1/a_n33_20# dff_10/dlatch_1/m1_27_49# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1079 m2_1376_n866# s2out dff_10/dlatch_1/nand_1/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1080 dff_10/dlatch_1/m1_27_49# clk vdd dff_10/dlatch_1/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1081 vdd dff_10/m1_n9_n58# dff_10/dlatch_1/m1_27_49# dff_10/dlatch_1/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1082 dff_10/dlatch_1/nand_0/a_n33_20# clk gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1083 dff_10/dlatch_1/m1_27_49# dff_10/m1_n9_n58# dff_10/dlatch_1/nand_0/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1084 dff_10/m1_n21_n58# dff_10/dlatch_0/m1_29_n71# vdd dff_10/dlatch_0/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1085 vdd dff_10/m1_n9_n58# dff_10/m1_n21_n58# dff_10/dlatch_0/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1086 dff_10/dlatch_0/nand_3/a_n33_20# dff_10/dlatch_0/m1_29_n71# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1087 dff_10/m1_n21_n58# dff_10/m1_n9_n58# dff_10/dlatch_0/nand_3/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1088 dff_10/dlatch_0/m1_29_n71# dff_10/m1_n65_174# vdd dff_10/dlatch_0/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1089 vdd s2 dff_10/dlatch_0/m1_29_n71# dff_10/dlatch_0/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1090 dff_10/dlatch_0/nand_2/a_n33_20# dff_10/m1_n65_174# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1091 dff_10/dlatch_0/m1_29_n71# s2 dff_10/dlatch_0/nand_2/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1092 dff_10/m1_n9_n58# dff_10/dlatch_0/m1_27_49# vdd dff_10/dlatch_0/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1093 vdd dff_10/m1_n21_n58# dff_10/m1_n9_n58# dff_10/dlatch_0/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1094 dff_10/dlatch_0/nand_1/a_n33_20# dff_10/dlatch_0/m1_27_49# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1095 dff_10/m1_n9_n58# dff_10/m1_n21_n58# dff_10/dlatch_0/nand_1/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1096 dff_10/dlatch_0/m1_27_49# dff_10/m1_n65_174# vdd dff_10/dlatch_0/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1097 vdd m1_1204_n278# dff_10/dlatch_0/m1_27_49# dff_10/dlatch_0/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1098 dff_10/dlatch_0/nand_0/a_n33_20# dff_10/m1_n65_174# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1099 dff_10/dlatch_0/m1_27_49# m1_1204_n278# dff_10/dlatch_0/nand_0/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1100 dff_10/m1_n65_174# clk vdd dff_10/inv_0/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1101 dff_10/m1_n65_174# clk gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1102 s1out dff_9/dlatch_1/m1_29_n71# vdd dff_9/dlatch_1/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1103 vdd m2_854_n873# s1out dff_9/dlatch_1/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1104 dff_9/dlatch_1/nand_3/a_n33_20# dff_9/dlatch_1/m1_29_n71# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1105 s1out m2_854_n873# dff_9/dlatch_1/nand_3/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1106 dff_9/dlatch_1/m1_29_n71# clk vdd dff_9/dlatch_1/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1107 vdd dff_9/m1_n21_n58# dff_9/dlatch_1/m1_29_n71# dff_9/dlatch_1/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1108 dff_9/dlatch_1/nand_2/a_n33_20# clk gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1109 dff_9/dlatch_1/m1_29_n71# dff_9/m1_n21_n58# dff_9/dlatch_1/nand_2/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1110 m2_854_n873# dff_9/dlatch_1/m1_27_49# vdd dff_9/dlatch_1/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1111 vdd s1out m2_854_n873# dff_9/dlatch_1/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1112 dff_9/dlatch_1/nand_1/a_n33_20# dff_9/dlatch_1/m1_27_49# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1113 m2_854_n873# s1out dff_9/dlatch_1/nand_1/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1114 dff_9/dlatch_1/m1_27_49# clk vdd dff_9/dlatch_1/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1115 vdd dff_9/m1_n9_n58# dff_9/dlatch_1/m1_27_49# dff_9/dlatch_1/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1116 dff_9/dlatch_1/nand_0/a_n33_20# clk gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1117 dff_9/dlatch_1/m1_27_49# dff_9/m1_n9_n58# dff_9/dlatch_1/nand_0/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1118 dff_9/m1_n21_n58# dff_9/dlatch_0/m1_29_n71# vdd dff_9/dlatch_0/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1119 vdd dff_9/m1_n9_n58# dff_9/m1_n21_n58# dff_9/dlatch_0/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1120 dff_9/dlatch_0/nand_3/a_n33_20# dff_9/dlatch_0/m1_29_n71# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1121 dff_9/m1_n21_n58# dff_9/m1_n9_n58# dff_9/dlatch_0/nand_3/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1122 dff_9/dlatch_0/m1_29_n71# dff_9/m1_n65_174# vdd dff_9/dlatch_0/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1123 vdd s1 dff_9/dlatch_0/m1_29_n71# dff_9/dlatch_0/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1124 dff_9/dlatch_0/nand_2/a_n33_20# dff_9/m1_n65_174# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1125 dff_9/dlatch_0/m1_29_n71# s1 dff_9/dlatch_0/nand_2/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1126 dff_9/m1_n9_n58# dff_9/dlatch_0/m1_27_49# vdd dff_9/dlatch_0/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1127 vdd dff_9/m1_n21_n58# dff_9/m1_n9_n58# dff_9/dlatch_0/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1128 dff_9/dlatch_0/nand_1/a_n33_20# dff_9/dlatch_0/m1_27_49# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1129 dff_9/m1_n9_n58# dff_9/m1_n21_n58# dff_9/dlatch_0/nand_1/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1130 dff_9/dlatch_0/m1_27_49# dff_9/m1_n65_174# vdd dff_9/dlatch_0/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1131 vdd m1_684_n288# dff_9/dlatch_0/m1_27_49# dff_9/dlatch_0/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1132 dff_9/dlatch_0/nand_0/a_n33_20# dff_9/m1_n65_174# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1133 dff_9/dlatch_0/m1_27_49# m1_684_n288# dff_9/dlatch_0/nand_0/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1134 dff_9/m1_n65_174# clk vdd dff_9/inv_0/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1135 dff_9/m1_n65_174# clk gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1136 cout dff_8/dlatch_1/m1_29_n71# vdd dff_8/dlatch_1/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1137 vdd m2_378_n882# cout dff_8/dlatch_1/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1138 dff_8/dlatch_1/nand_3/a_n33_20# dff_8/dlatch_1/m1_29_n71# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1139 cout m2_378_n882# dff_8/dlatch_1/nand_3/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1140 dff_8/dlatch_1/m1_29_n71# clk vdd dff_8/dlatch_1/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1141 vdd dff_8/m1_n21_n58# dff_8/dlatch_1/m1_29_n71# dff_8/dlatch_1/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1142 dff_8/dlatch_1/nand_2/a_n33_20# clk gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1143 dff_8/dlatch_1/m1_29_n71# dff_8/m1_n21_n58# dff_8/dlatch_1/nand_2/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1144 m2_378_n882# dff_8/dlatch_1/m1_27_49# vdd dff_8/dlatch_1/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1145 vdd cout m2_378_n882# dff_8/dlatch_1/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1146 dff_8/dlatch_1/nand_1/a_n33_20# dff_8/dlatch_1/m1_27_49# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1147 m2_378_n882# cout dff_8/dlatch_1/nand_1/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1148 dff_8/dlatch_1/m1_27_49# clk vdd dff_8/dlatch_1/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1149 vdd dff_8/m1_n9_n58# dff_8/dlatch_1/m1_27_49# dff_8/dlatch_1/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1150 dff_8/dlatch_1/nand_0/a_n33_20# clk gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1151 dff_8/dlatch_1/m1_27_49# dff_8/m1_n9_n58# dff_8/dlatch_1/nand_0/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1152 dff_8/m1_n21_n58# dff_8/dlatch_0/m1_29_n71# vdd dff_8/dlatch_0/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1153 vdd dff_8/m1_n9_n58# dff_8/m1_n21_n58# dff_8/dlatch_0/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1154 dff_8/dlatch_0/nand_3/a_n33_20# dff_8/dlatch_0/m1_29_n71# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1155 dff_8/m1_n21_n58# dff_8/m1_n9_n58# dff_8/dlatch_0/nand_3/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1156 dff_8/dlatch_0/m1_29_n71# dff_8/m1_n65_174# vdd dff_8/dlatch_0/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1157 vdd c4 dff_8/dlatch_0/m1_29_n71# dff_8/dlatch_0/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1158 dff_8/dlatch_0/nand_2/a_n33_20# dff_8/m1_n65_174# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1159 dff_8/dlatch_0/m1_29_n71# c4 dff_8/dlatch_0/nand_2/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1160 dff_8/m1_n9_n58# dff_8/dlatch_0/m1_27_49# vdd dff_8/dlatch_0/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1161 vdd dff_8/m1_n21_n58# dff_8/m1_n9_n58# dff_8/dlatch_0/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1162 dff_8/dlatch_0/nand_1/a_n33_20# dff_8/dlatch_0/m1_27_49# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1163 dff_8/m1_n9_n58# dff_8/m1_n21_n58# dff_8/dlatch_0/nand_1/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1164 dff_8/dlatch_0/m1_27_49# dff_8/m1_n65_174# vdd dff_8/dlatch_0/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1165 vdd m1_206_n285# dff_8/dlatch_0/m1_27_49# dff_8/dlatch_0/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1166 dff_8/dlatch_0/nand_0/a_n33_20# dff_8/m1_n65_174# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1167 dff_8/dlatch_0/m1_27_49# m1_206_n285# dff_8/dlatch_0/nand_0/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1168 dff_8/m1_n65_174# clk vdd dff_8/inv_0/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1169 dff_8/m1_n65_174# clk gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1170 m1_206_n285# c4 vdd inv_4/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1171 m1_206_n285# c4 m1_1815_211# Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=1200 ps=660
M1172 s4_inv s4 vdd inv_3/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1173 s4_inv s4 m1_1815_211# Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1174 m1_1732_n280# s3 vdd inv_2/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1175 m1_1732_n280# s3 m1_1815_211# Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1176 m1_1204_n278# s2 vdd inv_1/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1177 m1_1204_n278# s2 m1_1815_211# Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1178 m1_684_n288# s1 vdd inv_0/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1179 m1_684_n288# s1 m1_1815_211# Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1180 adder_0/lsum_0/xor_2/a_80_n16# adder_0/m1_846_n52# vdd adder_0/lsum_0/xor_2/inv_1/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1181 adder_0/lsum_0/xor_2/a_80_n16# adder_0/m1_846_n52# m1_1815_211# Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1182 adder_0/lsum_0/xor_2/a_72_n5# adder_0/m1_622_n582# vdd adder_0/lsum_0/xor_2/inv_0/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1183 adder_0/lsum_0/xor_2/a_72_n5# adder_0/m1_622_n582# m1_1815_211# Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1184 vdd adder_0/m1_622_n582# adder_0/lsum_0/xor_2/a_53_26# adder_0/lsum_0/xor_2/w_47_20# CMOSP w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M1185 adder_0/lsum_0/xor_2/a_53_26# adder_0/m1_846_n52# vdd adder_0/lsum_0/xor_2/w_47_20# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1186 s4 adder_0/lsum_0/xor_2/a_72_n5# adder_0/lsum_0/xor_2/a_53_26# adder_0/lsum_0/xor_2/w_47_20# CMOSP w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1187 adder_0/lsum_0/xor_2/a_53_26# adder_0/lsum_0/xor_2/a_80_n16# s4 adder_0/lsum_0/xor_2/w_47_20# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1188 adder_0/lsum_0/xor_2/a_60_n47# adder_0/m1_622_n582# m1_1815_211# Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1189 s4 adder_0/m1_846_n52# adder_0/lsum_0/xor_2/a_60_n47# Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1190 adder_0/lsum_0/xor_2/a_76_n47# adder_0/lsum_0/xor_2/a_72_n5# s4 Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1191 m1_1815_211# adder_0/lsum_0/xor_2/a_80_n16# adder_0/lsum_0/xor_2/a_76_n47# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1192 adder_0/lsum_0/xor_1/a_80_n16# adder_0/m1_684_n98# vdd adder_0/lsum_0/xor_1/inv_1/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1193 adder_0/lsum_0/xor_1/a_80_n16# adder_0/m1_684_n98# m1_1815_211# Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1194 adder_0/lsum_0/xor_1/a_72_n5# adder_0/m1_217_n553# vdd adder_0/lsum_0/xor_1/inv_0/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1195 adder_0/lsum_0/xor_1/a_72_n5# adder_0/m1_217_n553# m1_1815_211# Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1196 vdd adder_0/m1_217_n553# adder_0/lsum_0/xor_1/a_53_26# adder_0/lsum_0/xor_1/w_47_20# CMOSP w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M1197 adder_0/lsum_0/xor_1/a_53_26# adder_0/m1_684_n98# vdd adder_0/lsum_0/xor_1/w_47_20# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1198 s3 adder_0/lsum_0/xor_1/a_72_n5# adder_0/lsum_0/xor_1/a_53_26# adder_0/lsum_0/xor_1/w_47_20# CMOSP w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1199 adder_0/lsum_0/xor_1/a_53_26# adder_0/lsum_0/xor_1/a_80_n16# s3 adder_0/lsum_0/xor_1/w_47_20# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1200 adder_0/lsum_0/xor_1/a_60_n47# adder_0/m1_217_n553# m1_1815_211# Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1201 s3 adder_0/m1_684_n98# adder_0/lsum_0/xor_1/a_60_n47# Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1202 adder_0/lsum_0/xor_1/a_76_n47# adder_0/lsum_0/xor_1/a_72_n5# s3 Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1203 m1_1815_211# adder_0/lsum_0/xor_1/a_80_n16# adder_0/lsum_0/xor_1/a_76_n47# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1204 adder_0/lsum_0/xor_0/a_80_n16# adder_0/m1_519_n5# vdd adder_0/lsum_0/xor_0/inv_1/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1205 adder_0/lsum_0/xor_0/a_80_n16# adder_0/m1_519_n5# m1_1815_211# Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1206 adder_0/lsum_0/xor_0/a_72_n5# adder_0/m2_n46_n56# vdd adder_0/lsum_0/xor_0/inv_0/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1207 adder_0/lsum_0/xor_0/a_72_n5# adder_0/m2_n46_n56# m1_1815_211# Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1208 vdd adder_0/m2_n46_n56# adder_0/lsum_0/xor_0/a_53_26# adder_0/lsum_0/xor_0/w_47_20# CMOSP w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M1209 adder_0/lsum_0/xor_0/a_53_26# adder_0/m1_519_n5# vdd adder_0/lsum_0/xor_0/w_47_20# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1210 s2 adder_0/lsum_0/xor_0/a_72_n5# adder_0/lsum_0/xor_0/a_53_26# adder_0/lsum_0/xor_0/w_47_20# CMOSP w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1211 adder_0/lsum_0/xor_0/a_53_26# adder_0/lsum_0/xor_0/a_80_n16# s2 adder_0/lsum_0/xor_0/w_47_20# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1212 adder_0/lsum_0/xor_0/a_60_n47# adder_0/m2_n46_n56# m1_1815_211# Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1213 s2 adder_0/m1_519_n5# adder_0/lsum_0/xor_0/a_60_n47# Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1214 adder_0/lsum_0/xor_0/a_76_n47# adder_0/lsum_0/xor_0/a_72_n5# s2 Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1215 m1_1815_211# adder_0/lsum_0/xor_0/a_80_n16# adder_0/lsum_0/xor_0/a_76_n47# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1216 c4 adder_0/carry_0/or4_0/a_n41_8# vdd adder_0/carry_0/or4_0/inv_0/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1217 c4 adder_0/carry_0/or4_0/a_n41_8# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1218 adder_0/carry_0/or4_0/a_n41_60# m1_1815_211# vdd adder_0/carry_0/or4_0/w_n54_54# CMOSP w=80 l=2
+  ad=480 pd=172 as=0 ps=0
M1219 adder_0/carry_0/or4_0/a_n33_60# adder_0/carry_0/m1_843_59# adder_0/carry_0/or4_0/a_n41_60# adder_0/carry_0/or4_0/w_n54_54# CMOSP w=80 l=2
+  ad=480 pd=172 as=0 ps=0
M1220 adder_0/carry_0/or4_0/a_n25_60# adder_0/carry_0/m1_694_39# adder_0/carry_0/or4_0/a_n33_60# adder_0/carry_0/or4_0/w_n54_54# CMOSP w=80 l=2
+  ad=480 pd=172 as=0 ps=0
M1221 adder_0/carry_0/or4_0/a_n41_8# adder_0/m2_215_n71# adder_0/carry_0/or4_0/a_n25_60# adder_0/carry_0/or4_0/w_n54_54# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1222 adder_0/carry_0/or4_0/a_n41_8# m1_1815_211# gnd Gnd CMOSN w=10 l=2
+  ad=120 pd=64 as=0 ps=0
M1223 gnd adder_0/carry_0/m1_843_59# adder_0/carry_0/or4_0/a_n41_8# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1224 adder_0/carry_0/or4_0/a_n41_8# adder_0/carry_0/m1_694_39# gnd Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1225 gnd adder_0/m2_215_n71# adder_0/carry_0/or4_0/a_n41_8# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1226 adder_0/m1_622_n582# adder_0/carry_0/or3_0/a_n33_8# vdd adder_0/carry_0/or3_0/inv_0/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1227 adder_0/m1_622_n582# adder_0/carry_0/or3_0/a_n33_8# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1228 adder_0/carry_0/or3_0/a_n33_53# adder_0/carry_0/m1_361_n123# vdd adder_0/carry_0/or3_0/w_n46_47# CMOSP w=60 l=2
+  ad=360 pd=132 as=0 ps=0
M1229 adder_0/carry_0/or3_0/a_n25_53# adder_0/carry_0/m1_309_39# adder_0/carry_0/or3_0/a_n33_53# adder_0/carry_0/or3_0/w_n46_47# CMOSP w=60 l=2
+  ad=360 pd=132 as=0 ps=0
M1230 adder_0/carry_0/or3_0/a_n33_8# adder_0/m1_195_n109# adder_0/carry_0/or3_0/a_n25_53# adder_0/carry_0/or3_0/w_n46_47# CMOSP w=60 l=2
+  ad=300 pd=130 as=0 ps=0
M1231 adder_0/carry_0/or3_0/a_n33_8# adder_0/carry_0/m1_361_n123# gnd Gnd CMOSN w=10 l=2
+  ad=110 pd=62 as=0 ps=0
M1232 gnd adder_0/carry_0/m1_309_39# adder_0/carry_0/or3_0/a_n33_8# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1233 adder_0/carry_0/or3_0/a_n33_8# adder_0/m1_195_n109# gnd Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1234 adder_0/m1_217_n553# adder_0/carry_0/or2_0/a_n25_8# vdd adder_0/carry_0/or2_0/inv_0/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1235 adder_0/m1_217_n553# adder_0/carry_0/or2_0/a_n25_8# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1236 adder_0/carry_0/or2_0/a_n25_48# adder_0/carry_0/m1_n9_n92# vdd adder_0/carry_0/or2_0/w_n38_42# CMOSP w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1237 adder_0/carry_0/or2_0/a_n25_8# adder_0/m1_110_n137# adder_0/carry_0/or2_0/a_n25_48# adder_0/carry_0/or2_0/w_n38_42# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1238 adder_0/carry_0/or2_0/a_n25_8# adder_0/carry_0/m1_n9_n92# gnd Gnd CMOSN w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1239 gnd adder_0/m1_110_n137# adder_0/carry_0/or2_0/a_n25_8# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1240 m1_1815_211# adder_0/carry_0/and4_0/a_n41_32# vdd adder_0/carry_0/and4_0/inv_0/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1241 m1_1815_211# adder_0/carry_0/and4_0/a_n41_32# gnd Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1242 adder_0/carry_0/and4_0/a_n41_32# adder_0/m2_n46_n56# vdd adder_0/carry_0/and4_0/w_n54_26# CMOSP w=20 l=2
+  ad=240 pd=104 as=0 ps=0
M1243 vdd adder_0/m1_519_n5# adder_0/carry_0/and4_0/a_n41_32# adder_0/carry_0/and4_0/w_n54_26# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1244 adder_0/carry_0/and4_0/a_n41_32# adder_0/m1_684_n98# vdd adder_0/carry_0/and4_0/w_n54_26# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1245 vdd adder_0/m1_846_n52# adder_0/carry_0/and4_0/a_n41_32# adder_0/carry_0/and4_0/w_n54_26# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1246 adder_0/carry_0/and4_0/a_n41_n43# adder_0/m2_n46_n56# gnd Gnd CMOSN w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1247 adder_0/carry_0/and4_0/a_n33_n43# adder_0/m1_519_n5# adder_0/carry_0/and4_0/a_n41_n43# Gnd CMOSN w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1248 adder_0/carry_0/and4_0/a_n25_n43# adder_0/m1_684_n98# adder_0/carry_0/and4_0/a_n33_n43# Gnd CMOSN w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1249 adder_0/carry_0/and4_0/a_n41_32# adder_0/m1_846_n52# adder_0/carry_0/and4_0/a_n25_n43# Gnd CMOSN w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1250 adder_0/carry_0/m1_843_59# adder_0/carry_0/and3_1/a_n33_32# vdd adder_0/carry_0/and3_1/inv_0/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1251 adder_0/carry_0/m1_843_59# adder_0/carry_0/and3_1/a_n33_32# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1252 adder_0/carry_0/and3_1/a_n33_32# adder_0/m1_110_n137# vdd adder_0/carry_0/and3_1/w_n46_26# CMOSP w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M1253 vdd adder_0/m1_684_n98# adder_0/carry_0/and3_1/a_n33_32# adder_0/carry_0/and3_1/w_n46_26# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1254 adder_0/carry_0/and3_1/a_n33_32# adder_0/m1_846_n52# vdd adder_0/carry_0/and3_1/w_n46_26# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1255 adder_0/carry_0/and3_1/a_n33_n29# adder_0/m1_110_n137# gnd Gnd CMOSN w=31 l=2
+  ad=186 pd=74 as=0 ps=0
M1256 adder_0/carry_0/and3_1/a_n25_n29# adder_0/m1_684_n98# adder_0/carry_0/and3_1/a_n33_n29# Gnd CMOSN w=31 l=2
+  ad=186 pd=74 as=0 ps=0
M1257 adder_0/carry_0/and3_1/a_n33_32# adder_0/m1_846_n52# adder_0/carry_0/and3_1/a_n25_n29# Gnd CMOSN w=31 l=2
+  ad=155 pd=72 as=0 ps=0
M1258 adder_0/carry_0/m1_694_39# adder_0/carry_0/and2_2/a_n33_61# vdd adder_0/carry_0/and2_2/inv_0/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1259 adder_0/carry_0/m1_694_39# adder_0/carry_0/and2_2/a_n33_61# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1260 adder_0/carry_0/and2_2/a_n33_61# adder_0/m1_195_n109# vdd adder_0/carry_0/and2_2/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1261 vdd adder_0/m1_846_n52# adder_0/carry_0/and2_2/a_n33_61# adder_0/carry_0/and2_2/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1262 adder_0/carry_0/and2_2/a_n33_20# adder_0/m1_195_n109# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1263 adder_0/carry_0/and2_2/a_n33_61# adder_0/m1_846_n52# adder_0/carry_0/and2_2/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1264 adder_0/carry_0/m1_361_n123# adder_0/carry_0/and3_0/a_n33_32# vdd adder_0/carry_0/and3_0/inv_0/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1265 adder_0/carry_0/m1_361_n123# adder_0/carry_0/and3_0/a_n33_32# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1266 adder_0/carry_0/and3_0/a_n33_32# adder_0/m2_n46_n56# vdd adder_0/carry_0/and3_0/w_n46_26# CMOSP w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M1267 vdd adder_0/m1_519_n5# adder_0/carry_0/and3_0/a_n33_32# adder_0/carry_0/and3_0/w_n46_26# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1268 adder_0/carry_0/and3_0/a_n33_32# adder_0/m1_684_n98# vdd adder_0/carry_0/and3_0/w_n46_26# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1269 adder_0/carry_0/and3_0/a_n33_n29# adder_0/m2_n46_n56# gnd Gnd CMOSN w=31 l=2
+  ad=186 pd=74 as=0 ps=0
M1270 adder_0/carry_0/and3_0/a_n25_n29# adder_0/m1_519_n5# adder_0/carry_0/and3_0/a_n33_n29# Gnd CMOSN w=31 l=2
+  ad=186 pd=74 as=0 ps=0
M1271 adder_0/carry_0/and3_0/a_n33_32# adder_0/m1_684_n98# adder_0/carry_0/and3_0/a_n25_n29# Gnd CMOSN w=31 l=2
+  ad=155 pd=72 as=0 ps=0
M1272 adder_0/carry_0/m1_309_39# adder_0/carry_0/and2_1/a_n33_61# vdd adder_0/carry_0/and2_1/inv_0/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1273 adder_0/carry_0/m1_309_39# adder_0/carry_0/and2_1/a_n33_61# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1274 adder_0/carry_0/and2_1/a_n33_61# adder_0/m1_110_n137# vdd adder_0/carry_0/and2_1/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1275 vdd adder_0/m1_684_n98# adder_0/carry_0/and2_1/a_n33_61# adder_0/carry_0/and2_1/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1276 adder_0/carry_0/and2_1/a_n33_20# adder_0/m1_110_n137# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1277 adder_0/carry_0/and2_1/a_n33_61# adder_0/m1_684_n98# adder_0/carry_0/and2_1/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1278 adder_0/carry_0/m1_n9_n92# adder_0/carry_0/and2_0/a_n33_61# vdd adder_0/carry_0/and2_0/inv_0/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1279 adder_0/carry_0/m1_n9_n92# adder_0/carry_0/and2_0/a_n33_61# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1280 adder_0/carry_0/and2_0/a_n33_61# adder_0/m2_n46_n56# vdd adder_0/carry_0/and2_0/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1281 vdd adder_0/m1_519_n5# adder_0/carry_0/and2_0/a_n33_61# adder_0/carry_0/and2_0/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1282 adder_0/carry_0/and2_0/a_n33_20# adder_0/m2_n46_n56# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1283 adder_0/carry_0/and2_0/a_n33_61# adder_0/m1_519_n5# adder_0/carry_0/and2_0/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1284 adder_0/pg_0/xor_3/a_80_n16# a4 vdd adder_0/pg_0/xor_3/inv_1/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1285 adder_0/pg_0/xor_3/a_80_n16# a4 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1286 adder_0/pg_0/xor_3/a_72_n5# b4 vdd adder_0/pg_0/xor_3/inv_0/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1287 adder_0/pg_0/xor_3/a_72_n5# b4 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1288 vdd b4 adder_0/pg_0/xor_3/a_53_26# adder_0/pg_0/xor_3/w_47_20# CMOSP w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M1289 adder_0/pg_0/xor_3/a_53_26# a4 vdd adder_0/pg_0/xor_3/w_47_20# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1290 adder_0/m1_846_n52# adder_0/pg_0/xor_3/a_72_n5# adder_0/pg_0/xor_3/a_53_26# adder_0/pg_0/xor_3/w_47_20# CMOSP w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1291 adder_0/pg_0/xor_3/a_53_26# adder_0/pg_0/xor_3/a_80_n16# adder_0/m1_846_n52# adder_0/pg_0/xor_3/w_47_20# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1292 adder_0/pg_0/xor_3/a_60_n47# b4 gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1293 adder_0/m1_846_n52# a4 adder_0/pg_0/xor_3/a_60_n47# Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1294 adder_0/pg_0/xor_3/a_76_n47# adder_0/pg_0/xor_3/a_72_n5# adder_0/m1_846_n52# Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1295 gnd adder_0/pg_0/xor_3/a_80_n16# adder_0/pg_0/xor_3/a_76_n47# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1296 adder_0/pg_0/xor_2/a_80_n16# a3 vdd adder_0/pg_0/xor_2/inv_1/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1297 adder_0/pg_0/xor_2/a_80_n16# a3 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1298 adder_0/pg_0/xor_2/a_72_n5# b3 vdd adder_0/pg_0/xor_2/inv_0/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1299 adder_0/pg_0/xor_2/a_72_n5# b3 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1300 vdd b3 adder_0/pg_0/xor_2/a_53_26# adder_0/pg_0/xor_2/w_47_20# CMOSP w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M1301 adder_0/pg_0/xor_2/a_53_26# a3 vdd adder_0/pg_0/xor_2/w_47_20# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1302 adder_0/m1_684_n98# adder_0/pg_0/xor_2/a_72_n5# adder_0/pg_0/xor_2/a_53_26# adder_0/pg_0/xor_2/w_47_20# CMOSP w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1303 adder_0/pg_0/xor_2/a_53_26# adder_0/pg_0/xor_2/a_80_n16# adder_0/m1_684_n98# adder_0/pg_0/xor_2/w_47_20# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1304 adder_0/pg_0/xor_2/a_60_n47# b3 gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1305 adder_0/m1_684_n98# a3 adder_0/pg_0/xor_2/a_60_n47# Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1306 adder_0/pg_0/xor_2/a_76_n47# adder_0/pg_0/xor_2/a_72_n5# adder_0/m1_684_n98# Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1307 gnd adder_0/pg_0/xor_2/a_80_n16# adder_0/pg_0/xor_2/a_76_n47# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1308 adder_0/pg_0/xor_1/a_80_n16# a2 vdd adder_0/pg_0/xor_1/inv_1/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1309 adder_0/pg_0/xor_1/a_80_n16# a2 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1310 adder_0/pg_0/xor_1/a_72_n5# b2 vdd adder_0/pg_0/xor_1/inv_0/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1311 adder_0/pg_0/xor_1/a_72_n5# b2 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1312 vdd b2 adder_0/pg_0/xor_1/a_53_26# adder_0/pg_0/xor_1/w_47_20# CMOSP w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M1313 adder_0/pg_0/xor_1/a_53_26# a2 vdd adder_0/pg_0/xor_1/w_47_20# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1314 adder_0/m1_519_n5# adder_0/pg_0/xor_1/a_72_n5# adder_0/pg_0/xor_1/a_53_26# adder_0/pg_0/xor_1/w_47_20# CMOSP w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1315 adder_0/pg_0/xor_1/a_53_26# adder_0/pg_0/xor_1/a_80_n16# adder_0/m1_519_n5# adder_0/pg_0/xor_1/w_47_20# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1316 adder_0/pg_0/xor_1/a_60_n47# b2 gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1317 adder_0/m1_519_n5# a2 adder_0/pg_0/xor_1/a_60_n47# Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1318 adder_0/pg_0/xor_1/a_76_n47# adder_0/pg_0/xor_1/a_72_n5# adder_0/m1_519_n5# Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1319 gnd adder_0/pg_0/xor_1/a_80_n16# adder_0/pg_0/xor_1/a_76_n47# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1320 adder_0/pg_0/xor_0/a_80_n16# a1 vdd adder_0/pg_0/xor_0/inv_1/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1321 adder_0/pg_0/xor_0/a_80_n16# a1 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1322 adder_0/pg_0/xor_0/a_72_n5# b1 vdd adder_0/pg_0/xor_0/inv_0/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1323 adder_0/pg_0/xor_0/a_72_n5# b1 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1324 vdd b1 adder_0/pg_0/xor_0/a_53_26# adder_0/pg_0/xor_0/w_47_20# CMOSP w=40 l=2
+  ad=0 pd=0 as=640 ps=272
M1325 adder_0/pg_0/xor_0/a_53_26# a1 vdd adder_0/pg_0/xor_0/w_47_20# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1326 s1 adder_0/pg_0/xor_0/a_72_n5# adder_0/pg_0/xor_0/a_53_26# adder_0/pg_0/xor_0/w_47_20# CMOSP w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1327 adder_0/pg_0/xor_0/a_53_26# adder_0/pg_0/xor_0/a_80_n16# s1 adder_0/pg_0/xor_0/w_47_20# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1328 adder_0/pg_0/xor_0/a_60_n47# b1 gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1329 s1 a1 adder_0/pg_0/xor_0/a_60_n47# Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1330 adder_0/pg_0/xor_0/a_76_n47# adder_0/pg_0/xor_0/a_72_n5# s1 Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1331 gnd adder_0/pg_0/xor_0/a_80_n16# adder_0/pg_0/xor_0/a_76_n47# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1332 adder_0/m1_195_n109# adder_0/pg_0/and2_3/a_n33_61# vdd adder_0/pg_0/and2_3/inv_0/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1333 adder_0/m1_195_n109# adder_0/pg_0/and2_3/a_n33_61# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1334 adder_0/pg_0/and2_3/a_n33_61# b3 vdd adder_0/pg_0/and2_3/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1335 vdd a3 adder_0/pg_0/and2_3/a_n33_61# adder_0/pg_0/and2_3/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1336 adder_0/pg_0/and2_3/a_n33_20# b3 gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1337 adder_0/pg_0/and2_3/a_n33_61# a3 adder_0/pg_0/and2_3/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1338 adder_0/m2_n46_n56# adder_0/pg_0/and2_2/a_n33_61# vdd adder_0/pg_0/and2_2/inv_0/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1339 adder_0/m2_n46_n56# adder_0/pg_0/and2_2/a_n33_61# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1340 adder_0/pg_0/and2_2/a_n33_61# b1 vdd adder_0/pg_0/and2_2/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1341 vdd a1 adder_0/pg_0/and2_2/a_n33_61# adder_0/pg_0/and2_2/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1342 adder_0/pg_0/and2_2/a_n33_20# b1 gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1343 adder_0/pg_0/and2_2/a_n33_61# a1 adder_0/pg_0/and2_2/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1344 adder_0/m2_215_n71# adder_0/pg_0/and2_0/a_n33_61# vdd adder_0/pg_0/and2_0/inv_0/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1345 adder_0/m2_215_n71# adder_0/pg_0/and2_0/a_n33_61# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1346 adder_0/pg_0/and2_0/a_n33_61# b4 vdd adder_0/pg_0/and2_0/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1347 vdd a4 adder_0/pg_0/and2_0/a_n33_61# adder_0/pg_0/and2_0/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1348 adder_0/pg_0/and2_0/a_n33_20# b4 gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1349 adder_0/pg_0/and2_0/a_n33_61# a4 adder_0/pg_0/and2_0/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1350 adder_0/m1_110_n137# adder_0/pg_0/and2_1/a_n33_61# vdd adder_0/pg_0/and2_1/inv_0/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1351 adder_0/m1_110_n137# adder_0/pg_0/and2_1/a_n33_61# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1352 adder_0/pg_0/and2_1/a_n33_61# b2 vdd adder_0/pg_0/and2_1/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1353 vdd a2 adder_0/pg_0/and2_1/a_n33_61# adder_0/pg_0/and2_1/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1354 adder_0/pg_0/and2_1/a_n33_20# b2 gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1355 adder_0/pg_0/and2_1/a_n33_61# a2 adder_0/pg_0/and2_1/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1356 dff_7/dlatch_1/m1_70_41# dff_7/dlatch_1/m1_29_n71# vdd dff_7/dlatch_1/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1357 vdd b4 dff_7/dlatch_1/m1_70_41# dff_7/dlatch_1/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1358 dff_7/dlatch_1/nand_3/a_n33_20# dff_7/dlatch_1/m1_29_n71# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1359 dff_7/dlatch_1/m1_70_41# b4 dff_7/dlatch_1/nand_3/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1360 dff_7/dlatch_1/m1_29_n71# clk vdd dff_7/dlatch_1/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1361 vdd dff_7/m1_n21_n58# dff_7/dlatch_1/m1_29_n71# dff_7/dlatch_1/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1362 dff_7/dlatch_1/nand_2/a_n33_20# clk gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1363 dff_7/dlatch_1/m1_29_n71# dff_7/m1_n21_n58# dff_7/dlatch_1/nand_2/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1364 b4 dff_7/dlatch_1/m1_27_49# vdd dff_7/dlatch_1/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1365 vdd dff_7/dlatch_1/m1_70_41# b4 dff_7/dlatch_1/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1366 dff_7/dlatch_1/nand_1/a_n33_20# dff_7/dlatch_1/m1_27_49# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1367 b4 dff_7/dlatch_1/m1_70_41# dff_7/dlatch_1/nand_1/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1368 dff_7/dlatch_1/m1_27_49# clk vdd dff_7/dlatch_1/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1369 vdd dff_7/m1_n9_n58# dff_7/dlatch_1/m1_27_49# dff_7/dlatch_1/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1370 dff_7/dlatch_1/nand_0/a_n33_20# clk gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1371 dff_7/dlatch_1/m1_27_49# dff_7/m1_n9_n58# dff_7/dlatch_1/nand_0/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1372 dff_7/m1_n21_n58# dff_7/dlatch_0/m1_29_n71# vdd dff_7/dlatch_0/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1373 vdd dff_7/m1_n9_n58# dff_7/m1_n21_n58# dff_7/dlatch_0/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1374 dff_7/dlatch_0/nand_3/a_n33_20# dff_7/dlatch_0/m1_29_n71# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1375 dff_7/m1_n21_n58# dff_7/m1_n9_n58# dff_7/dlatch_0/nand_3/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1376 dff_7/dlatch_0/m1_29_n71# dff_7/m1_n65_174# vdd dff_7/dlatch_0/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1377 vdd b4in_inv dff_7/dlatch_0/m1_29_n71# dff_7/dlatch_0/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1378 dff_7/dlatch_0/nand_2/a_n33_20# dff_7/m1_n65_174# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1379 dff_7/dlatch_0/m1_29_n71# b4in_inv dff_7/dlatch_0/nand_2/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1380 dff_7/m1_n9_n58# dff_7/dlatch_0/m1_27_49# vdd dff_7/dlatch_0/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1381 vdd dff_7/m1_n21_n58# dff_7/m1_n9_n58# dff_7/dlatch_0/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1382 dff_7/dlatch_0/nand_1/a_n33_20# dff_7/dlatch_0/m1_27_49# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1383 dff_7/m1_n9_n58# dff_7/m1_n21_n58# dff_7/dlatch_0/nand_1/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1384 dff_7/dlatch_0/m1_27_49# dff_7/m1_n65_174# vdd dff_7/dlatch_0/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1385 vdd b4in dff_7/dlatch_0/m1_27_49# dff_7/dlatch_0/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1386 dff_7/dlatch_0/nand_0/a_n33_20# dff_7/m1_n65_174# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1387 dff_7/dlatch_0/m1_27_49# b4in dff_7/dlatch_0/nand_0/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1388 dff_7/m1_n65_174# clk vdd dff_7/inv_0/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1389 dff_7/m1_n65_174# clk gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1390 dff_6/dlatch_1/m1_70_41# dff_6/dlatch_1/m1_29_n71# vdd dff_6/dlatch_1/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1391 vdd a4 dff_6/dlatch_1/m1_70_41# dff_6/dlatch_1/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1392 dff_6/dlatch_1/nand_3/a_n33_20# dff_6/dlatch_1/m1_29_n71# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1393 dff_6/dlatch_1/m1_70_41# a4 dff_6/dlatch_1/nand_3/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1394 dff_6/dlatch_1/m1_29_n71# clk vdd dff_6/dlatch_1/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1395 vdd dff_6/m1_n21_n58# dff_6/dlatch_1/m1_29_n71# dff_6/dlatch_1/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1396 dff_6/dlatch_1/nand_2/a_n33_20# clk gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1397 dff_6/dlatch_1/m1_29_n71# dff_6/m1_n21_n58# dff_6/dlatch_1/nand_2/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1398 a4 dff_6/dlatch_1/m1_27_49# vdd dff_6/dlatch_1/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1399 vdd dff_6/dlatch_1/m1_70_41# a4 dff_6/dlatch_1/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1400 dff_6/dlatch_1/nand_1/a_n33_20# dff_6/dlatch_1/m1_27_49# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1401 a4 dff_6/dlatch_1/m1_70_41# dff_6/dlatch_1/nand_1/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1402 dff_6/dlatch_1/m1_27_49# clk vdd dff_6/dlatch_1/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1403 vdd dff_6/m1_n9_n58# dff_6/dlatch_1/m1_27_49# dff_6/dlatch_1/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1404 dff_6/dlatch_1/nand_0/a_n33_20# clk gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1405 dff_6/dlatch_1/m1_27_49# dff_6/m1_n9_n58# dff_6/dlatch_1/nand_0/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1406 dff_6/m1_n21_n58# dff_6/dlatch_0/m1_29_n71# vdd dff_6/dlatch_0/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1407 vdd dff_6/m1_n9_n58# dff_6/m1_n21_n58# dff_6/dlatch_0/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1408 dff_6/dlatch_0/nand_3/a_n33_20# dff_6/dlatch_0/m1_29_n71# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1409 dff_6/m1_n21_n58# dff_6/m1_n9_n58# dff_6/dlatch_0/nand_3/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1410 dff_6/dlatch_0/m1_29_n71# dff_6/m1_n65_174# vdd dff_6/dlatch_0/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1411 vdd a4in_inv dff_6/dlatch_0/m1_29_n71# dff_6/dlatch_0/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1412 dff_6/dlatch_0/nand_2/a_n33_20# dff_6/m1_n65_174# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1413 dff_6/dlatch_0/m1_29_n71# a4in_inv dff_6/dlatch_0/nand_2/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1414 dff_6/m1_n9_n58# dff_6/dlatch_0/m1_27_49# vdd dff_6/dlatch_0/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1415 vdd dff_6/m1_n21_n58# dff_6/m1_n9_n58# dff_6/dlatch_0/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1416 dff_6/dlatch_0/nand_1/a_n33_20# dff_6/dlatch_0/m1_27_49# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1417 dff_6/m1_n9_n58# dff_6/m1_n21_n58# dff_6/dlatch_0/nand_1/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1418 dff_6/dlatch_0/m1_27_49# dff_6/m1_n65_174# vdd dff_6/dlatch_0/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1419 vdd a4in dff_6/dlatch_0/m1_27_49# dff_6/dlatch_0/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1420 dff_6/dlatch_0/nand_0/a_n33_20# dff_6/m1_n65_174# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1421 dff_6/dlatch_0/m1_27_49# a4in dff_6/dlatch_0/nand_0/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1422 dff_6/m1_n65_174# clk vdd dff_6/inv_0/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1423 dff_6/m1_n65_174# clk gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1424 dff_5/dlatch_1/m1_70_41# dff_5/dlatch_1/m1_29_n71# vdd dff_5/dlatch_1/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1425 vdd b3 dff_5/dlatch_1/m1_70_41# dff_5/dlatch_1/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1426 dff_5/dlatch_1/nand_3/a_n33_20# dff_5/dlatch_1/m1_29_n71# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1427 dff_5/dlatch_1/m1_70_41# b3 dff_5/dlatch_1/nand_3/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1428 dff_5/dlatch_1/m1_29_n71# clk vdd dff_5/dlatch_1/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1429 vdd dff_5/m1_n21_n58# dff_5/dlatch_1/m1_29_n71# dff_5/dlatch_1/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1430 dff_5/dlatch_1/nand_2/a_n33_20# clk gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1431 dff_5/dlatch_1/m1_29_n71# dff_5/m1_n21_n58# dff_5/dlatch_1/nand_2/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1432 b3 dff_5/dlatch_1/m1_27_49# vdd dff_5/dlatch_1/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1433 vdd dff_5/dlatch_1/m1_70_41# b3 dff_5/dlatch_1/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1434 dff_5/dlatch_1/nand_1/a_n33_20# dff_5/dlatch_1/m1_27_49# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1435 b3 dff_5/dlatch_1/m1_70_41# dff_5/dlatch_1/nand_1/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1436 dff_5/dlatch_1/m1_27_49# clk vdd dff_5/dlatch_1/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1437 vdd dff_5/m1_n9_n58# dff_5/dlatch_1/m1_27_49# dff_5/dlatch_1/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1438 dff_5/dlatch_1/nand_0/a_n33_20# clk gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1439 dff_5/dlatch_1/m1_27_49# dff_5/m1_n9_n58# dff_5/dlatch_1/nand_0/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1440 dff_5/m1_n21_n58# dff_5/dlatch_0/m1_29_n71# vdd dff_5/dlatch_0/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1441 vdd dff_5/m1_n9_n58# dff_5/m1_n21_n58# dff_5/dlatch_0/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1442 dff_5/dlatch_0/nand_3/a_n33_20# dff_5/dlatch_0/m1_29_n71# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1443 dff_5/m1_n21_n58# dff_5/m1_n9_n58# dff_5/dlatch_0/nand_3/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1444 dff_5/dlatch_0/m1_29_n71# dff_5/m1_n65_174# vdd dff_5/dlatch_0/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1445 vdd b3in_inv dff_5/dlatch_0/m1_29_n71# dff_5/dlatch_0/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1446 dff_5/dlatch_0/nand_2/a_n33_20# dff_5/m1_n65_174# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1447 dff_5/dlatch_0/m1_29_n71# b3in_inv dff_5/dlatch_0/nand_2/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1448 dff_5/m1_n9_n58# dff_5/dlatch_0/m1_27_49# vdd dff_5/dlatch_0/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1449 vdd dff_5/m1_n21_n58# dff_5/m1_n9_n58# dff_5/dlatch_0/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1450 dff_5/dlatch_0/nand_1/a_n33_20# dff_5/dlatch_0/m1_27_49# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1451 dff_5/m1_n9_n58# dff_5/m1_n21_n58# dff_5/dlatch_0/nand_1/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1452 dff_5/dlatch_0/m1_27_49# dff_5/m1_n65_174# vdd dff_5/dlatch_0/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1453 vdd b3in dff_5/dlatch_0/m1_27_49# dff_5/dlatch_0/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1454 dff_5/dlatch_0/nand_0/a_n33_20# dff_5/m1_n65_174# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1455 dff_5/dlatch_0/m1_27_49# b3in dff_5/dlatch_0/nand_0/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1456 dff_5/m1_n65_174# clk vdd dff_5/inv_0/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1457 dff_5/m1_n65_174# clk gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1458 dff_4/dlatch_1/m1_70_41# dff_4/dlatch_1/m1_29_n71# vdd dff_4/dlatch_1/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1459 vdd a3 dff_4/dlatch_1/m1_70_41# dff_4/dlatch_1/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1460 dff_4/dlatch_1/nand_3/a_n33_20# dff_4/dlatch_1/m1_29_n71# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1461 dff_4/dlatch_1/m1_70_41# a3 dff_4/dlatch_1/nand_3/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1462 dff_4/dlatch_1/m1_29_n71# clk vdd dff_4/dlatch_1/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1463 vdd dff_4/m1_n21_n58# dff_4/dlatch_1/m1_29_n71# dff_4/dlatch_1/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1464 dff_4/dlatch_1/nand_2/a_n33_20# clk gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1465 dff_4/dlatch_1/m1_29_n71# dff_4/m1_n21_n58# dff_4/dlatch_1/nand_2/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1466 a3 dff_4/dlatch_1/m1_27_49# vdd dff_4/dlatch_1/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1467 vdd dff_4/dlatch_1/m1_70_41# a3 dff_4/dlatch_1/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1468 dff_4/dlatch_1/nand_1/a_n33_20# dff_4/dlatch_1/m1_27_49# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1469 a3 dff_4/dlatch_1/m1_70_41# dff_4/dlatch_1/nand_1/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1470 dff_4/dlatch_1/m1_27_49# clk vdd dff_4/dlatch_1/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1471 vdd dff_4/m1_n9_n58# dff_4/dlatch_1/m1_27_49# dff_4/dlatch_1/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1472 dff_4/dlatch_1/nand_0/a_n33_20# clk gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1473 dff_4/dlatch_1/m1_27_49# dff_4/m1_n9_n58# dff_4/dlatch_1/nand_0/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1474 dff_4/m1_n21_n58# dff_4/dlatch_0/m1_29_n71# vdd dff_4/dlatch_0/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1475 vdd dff_4/m1_n9_n58# dff_4/m1_n21_n58# dff_4/dlatch_0/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1476 dff_4/dlatch_0/nand_3/a_n33_20# dff_4/dlatch_0/m1_29_n71# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1477 dff_4/m1_n21_n58# dff_4/m1_n9_n58# dff_4/dlatch_0/nand_3/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1478 dff_4/dlatch_0/m1_29_n71# dff_4/m1_n65_174# vdd dff_4/dlatch_0/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1479 vdd a3in_inv dff_4/dlatch_0/m1_29_n71# dff_4/dlatch_0/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1480 dff_4/dlatch_0/nand_2/a_n33_20# dff_4/m1_n65_174# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1481 dff_4/dlatch_0/m1_29_n71# a3in_inv dff_4/dlatch_0/nand_2/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1482 dff_4/m1_n9_n58# dff_4/dlatch_0/m1_27_49# vdd dff_4/dlatch_0/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1483 vdd dff_4/m1_n21_n58# dff_4/m1_n9_n58# dff_4/dlatch_0/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1484 dff_4/dlatch_0/nand_1/a_n33_20# dff_4/dlatch_0/m1_27_49# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1485 dff_4/m1_n9_n58# dff_4/m1_n21_n58# dff_4/dlatch_0/nand_1/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1486 dff_4/dlatch_0/m1_27_49# dff_4/m1_n65_174# vdd dff_4/dlatch_0/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1487 vdd a3in dff_4/dlatch_0/m1_27_49# dff_4/dlatch_0/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1488 dff_4/dlatch_0/nand_0/a_n33_20# dff_4/m1_n65_174# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1489 dff_4/dlatch_0/m1_27_49# a3in dff_4/dlatch_0/nand_0/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1490 dff_4/m1_n65_174# clk vdd dff_4/inv_0/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1491 dff_4/m1_n65_174# clk gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1492 dff_3/dlatch_1/m1_70_41# dff_3/dlatch_1/m1_29_n71# vdd dff_3/dlatch_1/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1493 vdd b2 dff_3/dlatch_1/m1_70_41# dff_3/dlatch_1/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1494 dff_3/dlatch_1/nand_3/a_n33_20# dff_3/dlatch_1/m1_29_n71# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1495 dff_3/dlatch_1/m1_70_41# b2 dff_3/dlatch_1/nand_3/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1496 dff_3/dlatch_1/m1_29_n71# clk vdd dff_3/dlatch_1/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1497 vdd dff_3/m1_n21_n58# dff_3/dlatch_1/m1_29_n71# dff_3/dlatch_1/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1498 dff_3/dlatch_1/nand_2/a_n33_20# clk gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1499 dff_3/dlatch_1/m1_29_n71# dff_3/m1_n21_n58# dff_3/dlatch_1/nand_2/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1500 b2 dff_3/dlatch_1/m1_27_49# vdd dff_3/dlatch_1/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1501 vdd dff_3/dlatch_1/m1_70_41# b2 dff_3/dlatch_1/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1502 dff_3/dlatch_1/nand_1/a_n33_20# dff_3/dlatch_1/m1_27_49# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1503 b2 dff_3/dlatch_1/m1_70_41# dff_3/dlatch_1/nand_1/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1504 dff_3/dlatch_1/m1_27_49# clk vdd dff_3/dlatch_1/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1505 vdd dff_3/m1_n9_n58# dff_3/dlatch_1/m1_27_49# dff_3/dlatch_1/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1506 dff_3/dlatch_1/nand_0/a_n33_20# clk gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1507 dff_3/dlatch_1/m1_27_49# dff_3/m1_n9_n58# dff_3/dlatch_1/nand_0/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1508 dff_3/m1_n21_n58# dff_3/dlatch_0/m1_29_n71# vdd dff_3/dlatch_0/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1509 vdd dff_3/m1_n9_n58# dff_3/m1_n21_n58# dff_3/dlatch_0/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1510 dff_3/dlatch_0/nand_3/a_n33_20# dff_3/dlatch_0/m1_29_n71# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1511 dff_3/m1_n21_n58# dff_3/m1_n9_n58# dff_3/dlatch_0/nand_3/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1512 dff_3/dlatch_0/m1_29_n71# dff_3/m1_n65_174# vdd dff_3/dlatch_0/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1513 vdd b2in_inv dff_3/dlatch_0/m1_29_n71# dff_3/dlatch_0/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1514 dff_3/dlatch_0/nand_2/a_n33_20# dff_3/m1_n65_174# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1515 dff_3/dlatch_0/m1_29_n71# b2in_inv dff_3/dlatch_0/nand_2/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1516 dff_3/m1_n9_n58# dff_3/dlatch_0/m1_27_49# vdd dff_3/dlatch_0/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1517 vdd dff_3/m1_n21_n58# dff_3/m1_n9_n58# dff_3/dlatch_0/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1518 dff_3/dlatch_0/nand_1/a_n33_20# dff_3/dlatch_0/m1_27_49# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1519 dff_3/m1_n9_n58# dff_3/m1_n21_n58# dff_3/dlatch_0/nand_1/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1520 dff_3/dlatch_0/m1_27_49# dff_3/m1_n65_174# vdd dff_3/dlatch_0/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1521 vdd b2in dff_3/dlatch_0/m1_27_49# dff_3/dlatch_0/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1522 dff_3/dlatch_0/nand_0/a_n33_20# dff_3/m1_n65_174# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1523 dff_3/dlatch_0/m1_27_49# b2in dff_3/dlatch_0/nand_0/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1524 dff_3/m1_n65_174# clk vdd dff_3/inv_0/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1525 dff_3/m1_n65_174# clk gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1526 dff_2/dlatch_1/m1_70_41# dff_2/dlatch_1/m1_29_n71# vdd dff_2/dlatch_1/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1527 vdd a2 dff_2/dlatch_1/m1_70_41# dff_2/dlatch_1/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1528 dff_2/dlatch_1/nand_3/a_n33_20# dff_2/dlatch_1/m1_29_n71# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1529 dff_2/dlatch_1/m1_70_41# a2 dff_2/dlatch_1/nand_3/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1530 dff_2/dlatch_1/m1_29_n71# clk vdd dff_2/dlatch_1/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1531 vdd dff_2/m1_n21_n58# dff_2/dlatch_1/m1_29_n71# dff_2/dlatch_1/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1532 dff_2/dlatch_1/nand_2/a_n33_20# clk gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1533 dff_2/dlatch_1/m1_29_n71# dff_2/m1_n21_n58# dff_2/dlatch_1/nand_2/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1534 a2 dff_2/dlatch_1/m1_27_49# vdd dff_2/dlatch_1/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1535 vdd dff_2/dlatch_1/m1_70_41# a2 dff_2/dlatch_1/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1536 dff_2/dlatch_1/nand_1/a_n33_20# dff_2/dlatch_1/m1_27_49# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1537 a2 dff_2/dlatch_1/m1_70_41# dff_2/dlatch_1/nand_1/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1538 dff_2/dlatch_1/m1_27_49# clk vdd dff_2/dlatch_1/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1539 vdd dff_2/m1_n9_n58# dff_2/dlatch_1/m1_27_49# dff_2/dlatch_1/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1540 dff_2/dlatch_1/nand_0/a_n33_20# clk gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1541 dff_2/dlatch_1/m1_27_49# dff_2/m1_n9_n58# dff_2/dlatch_1/nand_0/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1542 dff_2/m1_n21_n58# dff_2/dlatch_0/m1_29_n71# vdd dff_2/dlatch_0/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1543 vdd dff_2/m1_n9_n58# dff_2/m1_n21_n58# dff_2/dlatch_0/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1544 dff_2/dlatch_0/nand_3/a_n33_20# dff_2/dlatch_0/m1_29_n71# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1545 dff_2/m1_n21_n58# dff_2/m1_n9_n58# dff_2/dlatch_0/nand_3/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1546 dff_2/dlatch_0/m1_29_n71# dff_2/m1_n65_174# vdd dff_2/dlatch_0/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1547 vdd a2in_inv dff_2/dlatch_0/m1_29_n71# dff_2/dlatch_0/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1548 dff_2/dlatch_0/nand_2/a_n33_20# dff_2/m1_n65_174# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1549 dff_2/dlatch_0/m1_29_n71# a2in_inv dff_2/dlatch_0/nand_2/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1550 dff_2/m1_n9_n58# dff_2/dlatch_0/m1_27_49# vdd dff_2/dlatch_0/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1551 vdd dff_2/m1_n21_n58# dff_2/m1_n9_n58# dff_2/dlatch_0/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1552 dff_2/dlatch_0/nand_1/a_n33_20# dff_2/dlatch_0/m1_27_49# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1553 dff_2/m1_n9_n58# dff_2/m1_n21_n58# dff_2/dlatch_0/nand_1/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1554 dff_2/dlatch_0/m1_27_49# dff_2/m1_n65_174# vdd dff_2/dlatch_0/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1555 vdd a2in dff_2/dlatch_0/m1_27_49# dff_2/dlatch_0/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1556 dff_2/dlatch_0/nand_0/a_n33_20# dff_2/m1_n65_174# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1557 dff_2/dlatch_0/m1_27_49# a2in dff_2/dlatch_0/nand_0/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1558 dff_2/m1_n65_174# clk vdd dff_2/inv_0/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1559 dff_2/m1_n65_174# clk gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1560 dff_1/dlatch_1/m1_70_41# dff_1/dlatch_1/m1_29_n71# vdd dff_1/dlatch_1/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1561 vdd b1 dff_1/dlatch_1/m1_70_41# dff_1/dlatch_1/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1562 dff_1/dlatch_1/nand_3/a_n33_20# dff_1/dlatch_1/m1_29_n71# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1563 dff_1/dlatch_1/m1_70_41# b1 dff_1/dlatch_1/nand_3/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1564 dff_1/dlatch_1/m1_29_n71# clk vdd dff_1/dlatch_1/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1565 vdd dff_1/m1_n21_n58# dff_1/dlatch_1/m1_29_n71# dff_1/dlatch_1/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1566 dff_1/dlatch_1/nand_2/a_n33_20# clk gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1567 dff_1/dlatch_1/m1_29_n71# dff_1/m1_n21_n58# dff_1/dlatch_1/nand_2/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1568 b1 dff_1/dlatch_1/m1_27_49# vdd dff_1/dlatch_1/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1569 vdd dff_1/dlatch_1/m1_70_41# b1 dff_1/dlatch_1/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1570 dff_1/dlatch_1/nand_1/a_n33_20# dff_1/dlatch_1/m1_27_49# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1571 b1 dff_1/dlatch_1/m1_70_41# dff_1/dlatch_1/nand_1/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1572 dff_1/dlatch_1/m1_27_49# clk vdd dff_1/dlatch_1/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1573 vdd dff_1/m1_n9_n58# dff_1/dlatch_1/m1_27_49# dff_1/dlatch_1/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1574 dff_1/dlatch_1/nand_0/a_n33_20# clk gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1575 dff_1/dlatch_1/m1_27_49# dff_1/m1_n9_n58# dff_1/dlatch_1/nand_0/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1576 dff_1/m1_n21_n58# dff_1/dlatch_0/m1_29_n71# vdd dff_1/dlatch_0/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1577 vdd dff_1/m1_n9_n58# dff_1/m1_n21_n58# dff_1/dlatch_0/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1578 dff_1/dlatch_0/nand_3/a_n33_20# dff_1/dlatch_0/m1_29_n71# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1579 dff_1/m1_n21_n58# dff_1/m1_n9_n58# dff_1/dlatch_0/nand_3/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1580 dff_1/dlatch_0/m1_29_n71# dff_1/m1_n65_174# vdd dff_1/dlatch_0/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1581 vdd b1in_inv dff_1/dlatch_0/m1_29_n71# dff_1/dlatch_0/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1582 dff_1/dlatch_0/nand_2/a_n33_20# dff_1/m1_n65_174# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1583 dff_1/dlatch_0/m1_29_n71# b1in_inv dff_1/dlatch_0/nand_2/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1584 dff_1/m1_n9_n58# dff_1/dlatch_0/m1_27_49# vdd dff_1/dlatch_0/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1585 vdd dff_1/m1_n21_n58# dff_1/m1_n9_n58# dff_1/dlatch_0/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1586 dff_1/dlatch_0/nand_1/a_n33_20# dff_1/dlatch_0/m1_27_49# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1587 dff_1/m1_n9_n58# dff_1/m1_n21_n58# dff_1/dlatch_0/nand_1/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1588 dff_1/dlatch_0/m1_27_49# dff_1/m1_n65_174# vdd dff_1/dlatch_0/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1589 vdd b1in dff_1/dlatch_0/m1_27_49# dff_1/dlatch_0/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1590 dff_1/dlatch_0/nand_0/a_n33_20# dff_1/m1_n65_174# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1591 dff_1/dlatch_0/m1_27_49# b1in dff_1/dlatch_0/nand_0/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1592 dff_1/m1_n65_174# clk vdd dff_1/inv_0/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1593 dff_1/m1_n65_174# clk gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1594 dff_0/dlatch_1/m1_70_41# dff_0/dlatch_1/m1_29_n71# vdd dff_0/dlatch_1/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1595 vdd a1 dff_0/dlatch_1/m1_70_41# dff_0/dlatch_1/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1596 dff_0/dlatch_1/nand_3/a_n33_20# dff_0/dlatch_1/m1_29_n71# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1597 dff_0/dlatch_1/m1_70_41# a1 dff_0/dlatch_1/nand_3/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1598 dff_0/dlatch_1/m1_29_n71# clk vdd dff_0/dlatch_1/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1599 vdd dff_0/m1_n21_n58# dff_0/dlatch_1/m1_29_n71# dff_0/dlatch_1/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1600 dff_0/dlatch_1/nand_2/a_n33_20# clk gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1601 dff_0/dlatch_1/m1_29_n71# dff_0/m1_n21_n58# dff_0/dlatch_1/nand_2/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1602 a1 dff_0/dlatch_1/m1_27_49# vdd dff_0/dlatch_1/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1603 vdd dff_0/dlatch_1/m1_70_41# a1 dff_0/dlatch_1/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1604 dff_0/dlatch_1/nand_1/a_n33_20# dff_0/dlatch_1/m1_27_49# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1605 a1 dff_0/dlatch_1/m1_70_41# dff_0/dlatch_1/nand_1/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1606 dff_0/dlatch_1/m1_27_49# clk vdd dff_0/dlatch_1/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1607 vdd dff_0/m1_n9_n58# dff_0/dlatch_1/m1_27_49# dff_0/dlatch_1/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1608 dff_0/dlatch_1/nand_0/a_n33_20# clk gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1609 dff_0/dlatch_1/m1_27_49# dff_0/m1_n9_n58# dff_0/dlatch_1/nand_0/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1610 dff_0/m1_n21_n58# dff_0/dlatch_0/m1_29_n71# vdd dff_0/dlatch_0/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1611 vdd dff_0/m1_n9_n58# dff_0/m1_n21_n58# dff_0/dlatch_0/nand_3/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1612 dff_0/dlatch_0/nand_3/a_n33_20# dff_0/dlatch_0/m1_29_n71# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1613 dff_0/m1_n21_n58# dff_0/m1_n9_n58# dff_0/dlatch_0/nand_3/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1614 dff_0/dlatch_0/m1_29_n71# dff_0/m1_n65_174# vdd dff_0/dlatch_0/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1615 vdd a1in_inv dff_0/dlatch_0/m1_29_n71# dff_0/dlatch_0/nand_2/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1616 dff_0/dlatch_0/nand_2/a_n33_20# dff_0/m1_n65_174# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1617 dff_0/dlatch_0/m1_29_n71# a1in_inv dff_0/dlatch_0/nand_2/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1618 dff_0/m1_n9_n58# dff_0/dlatch_0/m1_27_49# vdd dff_0/dlatch_0/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1619 vdd dff_0/m1_n21_n58# dff_0/m1_n9_n58# dff_0/dlatch_0/nand_1/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1620 dff_0/dlatch_0/nand_1/a_n33_20# dff_0/dlatch_0/m1_27_49# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1621 dff_0/m1_n9_n58# dff_0/m1_n21_n58# dff_0/dlatch_0/nand_1/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1622 dff_0/dlatch_0/m1_27_49# dff_0/m1_n65_174# vdd dff_0/dlatch_0/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1623 vdd a1in dff_0/dlatch_0/m1_27_49# dff_0/dlatch_0/nand_0/w_n46_55# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1624 dff_0/dlatch_0/nand_0/a_n33_20# dff_0/m1_n65_174# gnd Gnd CMOSN w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1625 dff_0/dlatch_0/m1_27_49# a1in dff_0/dlatch_0/nand_0/a_n33_20# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1626 dff_0/m1_n65_174# clk vdd dff_0/inv_0/w_n16_11# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1627 dff_0/m1_n65_174# clk gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
C0 adder_0/m1_217_n553# adder_0/m1_684_n98# 2.0fF
C1 b1 a1 4.7fF
C2 s4_inv s4 1.5fF
C3 vdd a3 1.5fF
C4 adder_0/m1_519_n5# adder_0/m1_684_n98# 3.2fF
C5 dff_12/m1_n21_n58# dff_12/m1_n9_n58# 1.3fF
C6 a4 vdd 1.1fF
C7 adder_0/m1_519_n5# adder_0/m1_110_n137# 1.0fF
C8 dff_9/m1_n21_n58# dff_9/m1_n9_n58# 1.3fF
C9 dff_4/m1_n21_n58# dff_4/m1_n9_n58# 1.3fF
C10 b2 a2 5.6fF
C11 vdd b2 1.0fF
C12 adder_0/carry_0/m1_843_59# adder_0/carry_0/m1_694_39# 1.5fF
C13 dff_7/m1_n21_n58# dff_7/m1_n9_n58# 1.3fF
C14 vdd a1 1.2fF
C15 c4 m1_206_n285# 4.2fF
C16 adder_0/m1_622_n582# adder_0/m1_846_n52# 1.9fF
C17 a4 b4 2.7fF
C18 m1_1204_n278# s2 1.1fF
C19 gnd vdd 2.7fF
C20 dff_0/m1_n21_n58# dff_0/m1_n9_n58# 1.3fF
C21 dff_11/m1_n21_n58# dff_11/m1_n9_n58# 1.3fF
C22 vdd b1 1.1fF
C23 dff_10/m1_n21_n58# dff_10/m1_n9_n58# 1.3fF
C24 vdd b3 1.2fF
C25 s3 s4 1.4fF
C26 adder_0/m1_846_n52# adder_0/m1_684_n98# 3.6fF
C27 dff_6/m1_n21_n58# dff_6/m1_n9_n58# 1.3fF
C28 m1_684_n288# s1 1.3fF
C29 vdd a2 1.0fF
C30 clk gnd 3.4fF
C31 adder_0/m1_684_n98# adder_0/m1_110_n137# 2.5fF
C32 adder_0/m1_684_n98# adder_0/m1_195_n109# 1.8fF
C33 adder_0/m2_n46_n56# vdd 1.6fF
C34 adder_0/m1_519_n5# adder_0/m2_n46_n56# 4.8fF
C35 b4 vdd 1.1fF
C36 adder_0/carry_0/m1_694_39# adder_0/m2_215_n71# 3.5fF
C37 dff_5/m1_n21_n58# dff_5/m1_n9_n58# 1.3fF
C38 dff_1/m1_n21_n58# dff_1/m1_n9_n58# 1.3fF
C39 dff_2/m1_n21_n58# dff_2/m1_n9_n58# 1.3fF
C40 adder_0/m1_195_n109# gnd 1.5fF
C41 clk vdd 2.9fF
C42 dff_8/m1_n21_n58# dff_8/m1_n9_n58# 1.3fF
C43 adder_0/carry_0/m1_309_39# adder_0/m1_195_n109# 1.4fF
C44 b3 a3 3.2fF
C45 a4 b3 7.0fF
C46 dff_3/m1_n21_n58# dff_3/m1_n9_n58# 1.3fF
C47 a1in gnd 2.0fF
C48 dff_0/m1_n65_174# gnd 2.6fF
C49 dff_0/dlatch_0/nand_0/w_n46_55# gnd 1.0fF
C50 dff_0/m1_n9_n58# gnd 6.1fF
C51 dff_0/m1_n21_n58# gnd 3.6fF
C52 dff_0/dlatch_0/nand_1/w_n46_55# gnd 1.0fF
C53 a1in_inv gnd 2.7fF
C54 dff_0/dlatch_0/nand_2/w_n46_55# gnd 1.0fF
C55 dff_0/dlatch_0/nand_3/w_n46_55# gnd 1.0fF
C56 dff_0/dlatch_1/nand_0/w_n46_55# gnd 1.0fF
C57 a1 gnd 13.8fF
C58 dff_0/dlatch_1/m1_70_41# gnd 1.3fF
C59 dff_0/dlatch_1/nand_1/w_n46_55# gnd 1.0fF
C60 dff_0/dlatch_1/nand_2/w_n46_55# gnd 1.0fF
C61 dff_0/dlatch_1/nand_3/w_n46_55# gnd 1.0fF
C62 b1in gnd 1.4fF
C63 dff_1/m1_n65_174# gnd 2.6fF
C64 dff_1/dlatch_0/nand_0/w_n46_55# gnd 1.0fF
C65 dff_1/m1_n9_n58# gnd 6.1fF
C66 dff_1/m1_n21_n58# gnd 3.6fF
C67 dff_1/dlatch_0/nand_1/w_n46_55# gnd 1.0fF
C68 b1in_inv gnd 5.1fF
C69 dff_1/dlatch_0/nand_2/w_n46_55# gnd 1.0fF
C70 dff_1/dlatch_0/nand_3/w_n46_55# gnd 1.0fF
C71 dff_1/dlatch_1/nand_0/w_n46_55# gnd 1.0fF
C72 b1 gnd 15.7fF
C73 dff_1/dlatch_1/m1_70_41# gnd 1.3fF
C74 dff_1/dlatch_1/nand_1/w_n46_55# gnd 1.0fF
C75 dff_1/dlatch_1/nand_2/w_n46_55# gnd 1.0fF
C76 dff_1/dlatch_1/nand_3/w_n46_55# gnd 1.0fF
C77 dff_2/m1_n65_174# gnd 2.6fF
C78 dff_2/dlatch_0/nand_0/w_n46_55# gnd 1.0fF
C79 dff_2/m1_n9_n58# gnd 6.1fF
C80 dff_2/m1_n21_n58# gnd 3.6fF
C81 dff_2/dlatch_0/nand_1/w_n46_55# gnd 1.0fF
C82 a2in_inv gnd 1.5fF
C83 dff_2/dlatch_0/nand_2/w_n46_55# gnd 1.0fF
C84 dff_2/dlatch_0/nand_3/w_n46_55# gnd 1.0fF
C85 dff_2/dlatch_1/nand_0/w_n46_55# gnd 1.0fF
C86 a2 gnd 19.3fF
C87 dff_2/dlatch_1/m1_70_41# gnd 1.3fF
C88 dff_2/dlatch_1/nand_1/w_n46_55# gnd 1.0fF
C89 dff_2/dlatch_1/nand_2/w_n46_55# gnd 1.0fF
C90 dff_2/dlatch_1/nand_3/w_n46_55# gnd 1.0fF
C91 dff_3/m1_n65_174# gnd 2.6fF
C92 dff_3/dlatch_0/nand_0/w_n46_55# gnd 1.0fF
C93 dff_3/m1_n9_n58# gnd 6.1fF
C94 dff_3/m1_n21_n58# gnd 3.6fF
C95 dff_3/dlatch_0/nand_1/w_n46_55# gnd 1.0fF
C96 b2in_inv gnd 1.6fF
C97 dff_3/dlatch_0/nand_2/w_n46_55# gnd 1.0fF
C98 dff_3/dlatch_0/nand_3/w_n46_55# gnd 1.0fF
C99 dff_3/dlatch_1/nand_0/w_n46_55# gnd 1.0fF
C100 b2 gnd 22.0fF
C101 dff_3/dlatch_1/m1_70_41# gnd 1.3fF
C102 dff_3/dlatch_1/nand_1/w_n46_55# gnd 1.0fF
C103 dff_3/dlatch_1/nand_2/w_n46_55# gnd 1.0fF
C104 dff_3/dlatch_1/nand_3/w_n46_55# gnd 1.0fF
C105 dff_4/m1_n65_174# gnd 2.6fF
C106 dff_4/dlatch_0/nand_0/w_n46_55# gnd 1.0fF
C107 dff_4/m1_n9_n58# gnd 6.1fF
C108 dff_4/m1_n21_n58# gnd 3.6fF
C109 dff_4/dlatch_0/nand_1/w_n46_55# gnd 1.0fF
C110 dff_4/dlatch_0/nand_2/w_n46_55# gnd 1.0fF
C111 dff_4/dlatch_0/nand_3/w_n46_55# gnd 1.0fF
C112 dff_4/dlatch_1/nand_0/w_n46_55# gnd 1.0fF
C113 a3 gnd 26.8fF
C114 dff_4/dlatch_1/m1_70_41# gnd 1.3fF
C115 dff_4/dlatch_1/nand_1/w_n46_55# gnd 1.0fF
C116 dff_4/dlatch_1/nand_2/w_n46_55# gnd 1.0fF
C117 dff_4/dlatch_1/nand_3/w_n46_55# gnd 1.0fF
C118 dff_5/m1_n65_174# gnd 2.6fF
C119 dff_5/dlatch_0/nand_0/w_n46_55# gnd 1.0fF
C120 dff_5/m1_n9_n58# gnd 6.1fF
C121 dff_5/m1_n21_n58# gnd 3.6fF
C122 dff_5/dlatch_0/nand_1/w_n46_55# gnd 1.0fF
C123 dff_5/dlatch_0/nand_2/w_n46_55# gnd 1.0fF
C124 dff_5/dlatch_0/nand_3/w_n46_55# gnd 1.0fF
C125 dff_5/dlatch_1/nand_0/w_n46_55# gnd 1.0fF
C126 b3 gnd 32.7fF
C127 dff_5/dlatch_1/m1_70_41# gnd 1.3fF
C128 dff_5/dlatch_1/nand_1/w_n46_55# gnd 1.0fF
C129 dff_5/dlatch_1/nand_2/w_n46_55# gnd 1.0fF
C130 dff_5/dlatch_1/nand_3/w_n46_55# gnd 1.0fF
C131 a4in gnd 7.6fF
C132 dff_6/m1_n65_174# gnd 2.6fF
C133 dff_6/dlatch_0/nand_0/w_n46_55# gnd 1.0fF
C134 dff_6/m1_n9_n58# gnd 6.1fF
C135 dff_6/m1_n21_n58# gnd 3.6fF
C136 dff_6/dlatch_0/nand_1/w_n46_55# gnd 1.0fF
C137 a4in_inv gnd 12.1fF
C138 dff_6/dlatch_0/nand_2/w_n46_55# gnd 1.0fF
C139 dff_6/dlatch_0/nand_3/w_n46_55# gnd 1.0fF
C140 dff_6/dlatch_1/nand_0/w_n46_55# gnd 1.0fF
C141 a4 gnd 34.0fF
C142 dff_6/dlatch_1/m1_70_41# gnd 1.3fF
C143 dff_6/dlatch_1/nand_1/w_n46_55# gnd 1.0fF
C144 dff_6/dlatch_1/nand_2/w_n46_55# gnd 1.0fF
C145 dff_6/dlatch_1/nand_3/w_n46_55# gnd 1.0fF
C146 b4in gnd 9.5fF
C147 dff_7/m1_n65_174# gnd 2.6fF
C148 dff_7/dlatch_0/nand_0/w_n46_55# gnd 1.0fF
C149 dff_7/m1_n9_n58# gnd 6.1fF
C150 dff_7/m1_n21_n58# gnd 3.6fF
C151 dff_7/dlatch_0/nand_1/w_n46_55# gnd 1.0fF
C152 b4in_inv gnd 14.7fF
C153 dff_7/dlatch_0/nand_2/w_n46_55# gnd 1.0fF
C154 dff_7/dlatch_0/nand_3/w_n46_55# gnd 1.0fF
C155 dff_7/dlatch_1/nand_0/w_n46_55# gnd 1.0fF
C156 dff_7/dlatch_1/m1_70_41# gnd 1.3fF
C157 dff_7/dlatch_1/nand_1/w_n46_55# gnd 1.0fF
C158 dff_7/dlatch_1/nand_2/w_n46_55# gnd 1.0fF
C159 dff_7/dlatch_1/nand_3/w_n46_55# gnd 1.0fF
C160 adder_0/pg_0/and2_1/w_n46_55# gnd 1.0fF
C161 adder_0/m1_110_n137# gnd 13.2fF
C162 adder_0/pg_0/and2_0/w_n46_55# gnd 1.0fF
C163 adder_0/m2_215_n71# gnd 12.9fF
C164 adder_0/pg_0/and2_2/w_n46_55# gnd 1.0fF
C165 adder_0/m2_n46_n56# gnd 42.1fF
C166 adder_0/pg_0/and2_3/w_n46_55# gnd 1.0fF
C167 adder_0/m1_195_n109# gnd 12.1fF
C168 adder_0/pg_0/xor_0/w_47_20# gnd 2.5fF
C169 adder_0/m1_519_n5# gnd 24.1fF
C170 adder_0/pg_0/xor_1/w_47_20# gnd 2.5fF
C171 adder_0/m1_684_n98# gnd 23.9fF
C172 adder_0/pg_0/xor_2/w_47_20# gnd 2.5fF
C173 adder_0/m1_846_n52# gnd 23.8fF
C174 adder_0/pg_0/xor_3/w_47_20# gnd 2.5fF
C175 adder_0/carry_0/and2_0/w_n46_55# gnd 1.0fF
C176 adder_0/carry_0/and2_1/w_n46_55# gnd 1.0fF
C177 adder_0/carry_0/m1_309_39# gnd 1.2fF
C178 adder_0/carry_0/and3_0/w_n46_26# gnd 1.3fF
C179 adder_0/carry_0/m1_361_n123# gnd 1.2fF
C180 adder_0/carry_0/and2_2/w_n46_55# gnd 1.0fF
C181 adder_0/carry_0/m1_694_39# gnd 1.6fF
C182 adder_0/carry_0/and3_1/w_n46_26# gnd 1.3fF
C183 adder_0/carry_0/m1_843_59# gnd 1.3fF
C184 adder_0/carry_0/and4_0/w_n54_26# gnd 1.5fF
C185 adder_0/carry_0/or2_0/w_n38_42# gnd 1.7fF
C186 adder_0/carry_0/or3_0/w_n46_47# gnd 2.9fF
C187 adder_0/carry_0/or4_0/w_n54_54# gnd 4.4fF
C188 adder_0/lsum_0/xor_0/w_47_20# gnd 2.5fF
C189 adder_0/lsum_0/xor_1/w_47_20# gnd 2.5fF
C190 adder_0/m1_217_n553# gnd 19.6fF
C191 adder_0/lsum_0/xor_2/w_47_20# gnd 2.5fF
C192 adder_0/m1_622_n582# gnd 16.1fF
C193 m1_684_n288# gnd 19.9fF
C194 s1 gnd 14.3fF
C195 m1_1204_n278# gnd 17.0fF
C196 s2 gnd 16.1fF
C197 m1_1732_n280# gnd 11.0fF
C198 s3 gnd 15.6fF
C199 s4_inv gnd 14.0fF
C200 s4 gnd 25.0fF
C201 m1_1815_211# gnd 9.4fF
C202 m1_206_n285# gnd 20.1fF
C203 c4 gnd 30.9fF
C204 dff_8/m1_n65_174# gnd 2.6fF
C205 dff_8/dlatch_0/nand_0/w_n46_55# gnd 1.0fF
C206 dff_8/m1_n9_n58# gnd 6.1fF
C207 dff_8/m1_n21_n58# gnd 3.6fF
C208 dff_8/dlatch_0/nand_1/w_n46_55# gnd 1.0fF
C209 dff_8/dlatch_0/nand_2/w_n46_55# gnd 1.0fF
C210 dff_8/dlatch_0/nand_3/w_n46_55# gnd 1.0fF
C211 dff_8/dlatch_1/nand_0/w_n46_55# gnd 1.0fF
C212 m2_378_n882# gnd 4.9fF
C213 cout gnd 2.0fF
C214 dff_8/dlatch_1/nand_1/w_n46_55# gnd 1.0fF
C215 dff_8/dlatch_1/nand_2/w_n46_55# gnd 1.0fF
C216 dff_8/dlatch_1/nand_3/w_n46_55# gnd 1.0fF
C217 dff_9/m1_n65_174# gnd 2.6fF
C218 dff_9/dlatch_0/nand_0/w_n46_55# gnd 1.0fF
C219 dff_9/m1_n9_n58# gnd 6.1fF
C220 dff_9/m1_n21_n58# gnd 3.6fF
C221 dff_9/dlatch_0/nand_1/w_n46_55# gnd 1.0fF
C222 dff_9/dlatch_0/nand_2/w_n46_55# gnd 1.0fF
C223 dff_9/dlatch_0/nand_3/w_n46_55# gnd 1.0fF
C224 dff_9/dlatch_1/nand_0/w_n46_55# gnd 1.0fF
C225 m2_854_n873# gnd 4.7fF
C226 s1out gnd 1.9fF
C227 dff_9/dlatch_1/nand_1/w_n46_55# gnd 1.0fF
C228 dff_9/dlatch_1/nand_2/w_n46_55# gnd 1.0fF
C229 dff_9/dlatch_1/nand_3/w_n46_55# gnd 1.0fF
C230 dff_10/m1_n65_174# gnd 2.6fF
C231 dff_10/dlatch_0/nand_0/w_n46_55# gnd 1.0fF
C232 dff_10/m1_n9_n58# gnd 6.1fF
C233 dff_10/m1_n21_n58# gnd 3.6fF
C234 dff_10/dlatch_0/nand_1/w_n46_55# gnd 1.0fF
C235 dff_10/dlatch_0/nand_2/w_n46_55# gnd 1.0fF
C236 dff_10/dlatch_0/nand_3/w_n46_55# gnd 1.0fF
C237 dff_10/dlatch_1/nand_0/w_n46_55# gnd 1.0fF
C238 m2_1376_n866# gnd 4.8fF
C239 s2out gnd 1.9fF
C240 dff_10/dlatch_1/nand_1/w_n46_55# gnd 1.0fF
C241 dff_10/dlatch_1/nand_2/w_n46_55# gnd 1.0fF
C242 dff_10/dlatch_1/nand_3/w_n46_55# gnd 1.0fF
C243 dff_11/m1_n65_174# gnd 2.6fF
C244 dff_11/dlatch_0/nand_0/w_n46_55# gnd 1.0fF
C245 dff_11/m1_n9_n58# gnd 6.1fF
C246 dff_11/m1_n21_n58# gnd 3.6fF
C247 dff_11/dlatch_0/nand_1/w_n46_55# gnd 1.0fF
C248 dff_11/dlatch_0/nand_2/w_n46_55# gnd 1.0fF
C249 dff_11/dlatch_0/nand_3/w_n46_55# gnd 1.0fF
C250 dff_11/dlatch_1/nand_0/w_n46_55# gnd 1.0fF
C251 m2_1903_n872# gnd 4.8fF
C252 s3out gnd 1.8fF
C253 dff_11/dlatch_1/nand_1/w_n46_55# gnd 1.0fF
C254 dff_11/dlatch_1/nand_2/w_n46_55# gnd 1.0fF
C255 dff_11/dlatch_1/nand_3/w_n46_55# gnd 1.0fF
C256 dff_12/m1_n65_174# gnd 2.6fF
C257 dff_12/dlatch_0/nand_0/w_n46_55# gnd 1.0fF
C258 dff_12/m1_n9_n58# gnd 6.1fF
C259 dff_12/m1_n21_n58# gnd 3.6fF
C260 dff_12/dlatch_0/nand_1/w_n46_55# gnd 1.0fF
C261 dff_12/dlatch_0/nand_2/w_n46_55# gnd 1.0fF
C262 dff_12/dlatch_0/nand_3/w_n46_55# gnd 1.0fF
C263 dff_12/dlatch_1/nand_0/w_n46_55# gnd 1.0fF
C264 m2_2425_n861# gnd 4.8fF
C265 s4out gnd 1.7fF
.ic v(clk) = 0
.tran 0.1ns 180n
.control
set hcopypscolor = 1
set color0=white
set color1=black

run
plot v(clk)
plot v(a4in)+6 v(a3in)+4 v(a2in)+2 v(a1in)
plot v(b4in)+6 v(b3in)+4 v(b2in)+2 v(b1in)
plot v(cout)+8 v(s4out)+6 v(s3out)+4 v(s2out)+2 v(s1out)
plot v(c4)+8 v(s4)+6 v(s3)+4 v(s2)+2 v(s1)
plot v(a4)+6 v(a3)+4 v(a2)+2 v(a1)
plot v(b4)+6 v(b3)+4 v(b2)+2 v(b1)
set curplottitle= "Aravind Narayanan-2019102014"

.endc
