magic
tech scmos
timestamp 1619483019
<< nwell >>
rect -1 0 101 39
<< ntransistor >>
rect 10 -32 12 -22
rect 27 -32 29 -22
rect 45 -32 47 -22
rect 64 -32 66 -22
rect 71 -32 73 -22
rect 88 -32 90 -22
<< ptransistor >>
rect 10 6 12 26
rect 28 6 30 26
rect 38 6 40 26
rect 64 6 66 26
rect 71 6 73 26
rect 88 6 90 26
<< ndiffusion >>
rect 9 -32 10 -22
rect 12 -32 13 -22
rect 26 -32 27 -22
rect 29 -32 45 -22
rect 47 -32 50 -22
rect 63 -32 64 -22
rect 66 -32 71 -22
rect 73 -32 74 -22
rect 87 -32 88 -22
rect 90 -32 91 -22
<< pdiffusion >>
rect 9 6 10 26
rect 12 6 13 26
rect 27 6 28 26
rect 30 6 38 26
rect 40 6 41 26
rect 63 6 64 26
rect 66 6 71 26
rect 73 6 74 26
rect 87 6 88 26
rect 90 6 91 26
<< ndcontact >>
rect 5 -32 9 -22
rect 13 -32 17 -22
rect 22 -32 26 -22
rect 50 -32 54 -22
rect 58 -32 63 -22
rect 74 -32 78 -22
rect 83 -32 87 -22
rect 91 -32 95 -22
<< pdcontact >>
rect 5 6 9 26
rect 13 6 17 26
rect 23 6 27 26
rect 41 6 45 26
rect 58 6 63 26
rect 74 6 78 26
rect 83 6 87 26
rect 91 6 95 26
<< polysilicon >>
rect 38 32 90 34
rect 10 26 12 29
rect 28 26 30 29
rect 38 26 40 32
rect 64 26 66 29
rect 71 26 73 29
rect 88 26 90 32
rect 10 -22 12 6
rect 28 -14 30 6
rect 38 5 40 6
rect 18 -16 30 -14
rect 37 3 40 5
rect 10 -35 12 -32
rect 18 -38 20 -16
rect 37 -19 39 3
rect 64 -10 66 6
rect 47 -12 66 -10
rect 27 -21 39 -19
rect 27 -22 29 -21
rect 45 -22 47 -12
rect 64 -22 66 -19
rect 71 -22 73 6
rect 88 -17 90 6
rect 88 -19 94 -17
rect 88 -22 90 -19
rect 27 -35 29 -32
rect 45 -35 47 -32
rect 64 -38 66 -32
rect 71 -35 73 -32
rect 88 -35 90 -32
rect 18 -40 66 -38
<< polycontact >>
rect 6 -5 10 -1
rect 24 -5 28 -1
rect 43 -12 47 -8
rect 73 -17 77 -12
rect 94 -19 98 -15
<< metal1 >>
rect -1 36 101 39
rect 5 26 9 36
rect 23 26 27 36
rect 74 26 78 36
rect 91 26 95 36
rect 13 -1 17 6
rect 41 -1 45 6
rect 58 -1 63 6
rect -1 -5 6 -1
rect 13 -5 24 -1
rect 41 -5 58 -1
rect 0 -7 5 -5
rect 13 -22 17 -5
rect 50 -6 58 -5
rect 50 -22 54 -6
rect 58 -22 63 -6
rect 83 -12 87 6
rect 77 -17 87 -12
rect 83 -22 87 -17
rect 5 -42 9 -32
rect 22 -42 26 -32
rect 74 -42 78 -32
rect 91 -42 95 -32
rect -1 -45 101 -42
<< m2contact >>
rect 0 -12 5 -7
rect 58 -6 63 -1
<< metal2 >>
rect 63 -6 101 -1
rect 5 -12 47 -8
<< labels >>
rlabel metal1 1 -4 1 -4 3 A
rlabel metal1 51 -44 51 -44 1 gnd
rlabel metal2 97 -4 97 -4 7 out
rlabel metal1 54 37 54 37 5 vdd
rlabel metal1 84 -15 84 -15 1 b_bar
rlabel metal1 16 -3 16 -3 1 a_bar
rlabel polycontact 96 -17 96 -17 7 B
<< end >>
