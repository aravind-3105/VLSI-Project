magic
tech scmos
timestamp 1619593969
<< nwell >>
rect 0 -1 34 51
<< ntransistor >>
rect 11 -35 13 -25
rect 19 -35 21 -25
<< ptransistor >>
rect 11 5 13 45
rect 19 5 21 45
<< ndiffusion >>
rect 10 -35 11 -25
rect 13 -35 14 -25
rect 18 -35 19 -25
rect 21 -35 22 -25
<< pdiffusion >>
rect 10 5 11 45
rect 13 5 19 45
rect 21 5 24 45
<< ndcontact >>
rect 6 -35 10 -25
rect 14 -35 18 -25
rect 22 -35 26 -25
<< pdcontact >>
rect 6 5 10 45
rect 24 5 28 45
<< polysilicon >>
rect 11 45 13 48
rect 19 45 21 48
rect 11 -11 13 5
rect 19 -4 21 5
rect 11 -25 13 -15
rect 19 -25 21 -8
rect 11 -38 13 -35
rect 19 -38 21 -35
<< polycontact >>
rect 17 -8 21 -4
rect 9 -15 13 -11
<< metal1 >>
rect 0 49 34 52
rect 6 45 10 49
rect 0 -8 17 -4
rect 24 -9 28 5
rect 0 -15 9 -11
rect 24 -13 34 -9
rect 24 -18 28 -13
rect 14 -22 28 -18
rect 14 -25 18 -22
rect 6 -39 10 -35
rect 22 -39 26 -35
rect -1 -42 34 -39
<< end >>
