.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.param W = {10*LAMBDA}
.param width_N={10*LAMBDA}
.param width_P={20*LAMBDA}
.global gnd vdd

Vdd	vdd	gnd	'SUPPLY'
vd10     P1     0 pulse 1.8 0 0ns  100ps 100ps 20ns  40ns
vd20     G1     0 pulse 1.8 0 0ns  100ps 100ps 30ns  40ns
vd11     P2     0 pulse 0 1.8 10ns 100ps 100ps 10ns  40ns
vd21     G2     0 pulse 1.8 0 0ns 100ps 100ps 30ns  40ns
vd12     P3     0 pulse 1.8 0 0ns 100ps 100ps 50ns  60ns
vd22     G3     0 pulse 1.8 0 0ns 100ps 100ps 20ns  30ns
vd13     P4     0 pulse 1.8 0 0ns 100ps 100ps 20ns  30ns
vd23     G4     0 pulse 1.8 0 0ns 100ps 100ps 40ns  60ns

vdC Ci 0 pulse 0 0 0ns 100ps 100ps 20ns 60ns

.subckt xor_subckt a b y vdd gnd
//Top inverter
M1      a_bar       a       vdd     vdd  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
M2      a_bar       a       gnd     gnd  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

//Bottom Inverter
M3      b_bar       b       vdd     vdd  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
M4      b_bar       b       gnd     gnd  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

//Layer 2
M5      J1   a_bar    vdd     vdd  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
M6      y       b       J1     J1  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
M7      y       a       J2     J2  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
M8      J2      b     gnd     gnd  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

//Layer 3
M9      J11       b_bar    vdd     vdd  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
M10      y       a         J11     J11  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
M11      y     a_bar       J22     J22  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
M12      J22     b_bar     gnd     gnd  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
.ends xor_subckt


.subckt and_subckt a b y vdd gnd
.param w_AND_P = {2*W}
.param w_AND_N = {2*W}
* Layer-1
M1      nand       b       vdd     vdd  CMOSP   W={w_AND_P}   L={2*LAMBDA}
+ AS={5*w_AND_P*LAMBDA} PS={10*LAMBDA+2*w_AND_P} AD={5*w_AND_P*LAMBDA} PD={10*LAMBDA+2*w_AND_P}
M2      nand       a       vdd     vdd  CMOSP   W={w_AND_P}   L={2*LAMBDA}
+ AS={5*w_AND_P*LAMBDA} PS={10*LAMBDA+2*w_AND_P} AD={5*w_AND_P*LAMBDA} PD={10*LAMBDA+2*w_AND_P}
M3      nand       a       J     J  CMOSN   W={w_AND_N}   L={2*LAMBDA}
+ AS={5*w_AND_N*LAMBDA} PS={10*LAMBDA+2*w_AND_N} AD={5*w_AND_N*LAMBDA} PD={10*LAMBDA+2*w_AND_N}
M4      J         b      gnd gnd   CMOSN   W={w_AND_N}   L={2*LAMBDA}
+ AS={5*w_AND_N*LAMBDA} PS={10*LAMBDA+2*w_AND_N} AD={5*w_AND_N*LAMBDA} PD={10*LAMBDA+2*w_AND_N}

M5      y       nand       vdd     vdd  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
M6      y       nand       gnd     gnd  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
.ends and_subckt

.subckt or_subckt a b y vdd gnd
.param w_OR_P = {4*W}
.param w_OR_N = {W}
* Layer-1
M1      J1       a       vdd     vdd  CMOSP   W={w_OR_P}   L={2*LAMBDA}
+ AS={5*w_OR_P*LAMBDA} PS={10*LAMBDA+2*w_OR_P} AD={5*w_OR_P*LAMBDA} PD={10*LAMBDA+2*w_OR_P}
M2      nor      b       J1      J1  CMOSP   W={w_OR_P}   L={2*LAMBDA}
+ AS={5*w_OR_P*LAMBDA} PS={10*LAMBDA+2*w_OR_P} AD={5*w_OR_P*LAMBDA} PD={10*LAMBDA+2*w_OR_P}
M3      nor       a     gnd   gnd   CMOSN   W={w_OR_N}   L={2*LAMBDA}
+ AS={5*w_OR_N*LAMBDA} PS={10*LAMBDA+2*w_OR_N} AD={5*w_OR_N*LAMBDA} PD={10*LAMBDA+2*w_OR_N}
M4      nor       b     gnd   gnd   CMOSN   W={w_OR_N}   L={2*LAMBDA}
+ AS={5*w_OR_N*LAMBDA} PS={10*LAMBDA+2*w_OR_N} AD={5*w_OR_N*LAMBDA} PD={10*LAMBDA+2*w_OR_N}

M5      y       nor       vdd     vdd  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
M6      y       nor       gnd     gnd  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
.ends or_subckt

.subckt or3_subckt a b c y vdd gnd
.param w_OR_P3 = {6*W}
.param w_OR_N3 = {W}
// NOR
M1      J1       a       vdd     vdd  CMOSP   W={w_OR_P3}   L={2*LAMBDA}
+ AS={5*w_OR_P3*LAMBDA} PS={10*LAMBDA+2*w_OR_P3} AD={5*w_OR_P3*LAMBDA} PD={10*LAMBDA+2*w_OR_P3}

M2      J2       b       J1      J1  CMOSP   W={w_OR_P3}   L={2*LAMBDA}
+ AS={5*w_OR_P3*LAMBDA} PS={10*LAMBDA+2*w_OR_P3} AD={5*w_OR_P3*LAMBDA} PD={10*LAMBDA+2*w_OR_P3}

M3      nor      c       J2      J2  CMOSP   W={w_OR_P3}   L={2*LAMBDA}
+ AS={5*w_OR_P3*LAMBDA} PS={10*LAMBDA+2*w_OR_P3} AD={5*w_OR_P3*LAMBDA} PD={10*LAMBDA+2*w_OR_P3}

M4      nor       a     gnd   gnd   CMOSN   W={w_OR_N3}   L={2*LAMBDA}
+ AS={5*w_OR_N3*LAMBDA} PS={10*LAMBDA+2*w_OR_N3} AD={5*w_OR_N3*LAMBDA} PD={10*LAMBDA+2*w_OR_N3}

M5      nor       b     gnd   gnd   CMOSN   W={w_OR_N3}   L={2*LAMBDA}
+ AS={5*w_OR_N3*LAMBDA} PS={10*LAMBDA+2*w_OR_N3} AD={5*w_OR_N3*LAMBDA} PD={10*LAMBDA+2*w_OR_N3}

M6      nor       c     gnd   gnd   CMOSN   W={w_OR_N3}   L={2*LAMBDA}
+ AS={5*w_OR_N3*LAMBDA} PS={10*LAMBDA+2*w_OR_N3} AD={5*w_OR_N3*LAMBDA} PD={10*LAMBDA+2*w_OR_N3}

// Inverter
M7      y       nor       vdd     vdd  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

M8      y       nor       gnd     gnd  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
.ends or3_subckt

.subckt or4_subckt a b c d y vdd gnd
.param w_OR_P4 = {8*W}
.param w_OR_N4 = {W}
// NOR
M1      J1       a       vdd     vdd  CMOSP   W={w_OR_P4}   L={2*LAMBDA}
+ AS={5*w_OR_P4*LAMBDA} PS={10*LAMBDA+2*w_OR_P4} AD={5*w_OR_P4*LAMBDA} PD={10*LAMBDA+2*w_OR_P4}

M2      J2       b       J1      J1  CMOSP   W={w_OR_P4}   L={2*LAMBDA}
+ AS={5*w_OR_P4*LAMBDA} PS={10*LAMBDA+2*w_OR_P4} AD={5*w_OR_P4*LAMBDA} PD={10*LAMBDA+2*w_OR_P4}

M3      J3       c       J2      J2  CMOSP   W={w_OR_P4}   L={2*LAMBDA}
+ AS={5*w_OR_P4*LAMBDA} PS={10*LAMBDA+2*w_OR_P4} AD={5*w_OR_P4*LAMBDA} PD={10*LAMBDA+2*w_OR_P4}

M4      nor      d       J3      J3  CMOSP   W={w_OR_P4}   L={2*LAMBDA}
+ AS={5*w_OR_P4*LAMBDA} PS={10*LAMBDA+2*w_OR_P4} AD={5*w_OR_P4*LAMBDA} PD={10*LAMBDA+2*w_OR_P4}

M5      nor       a     gnd   gnd   CMOSN   W={w_OR_N4}   L={2*LAMBDA}
+ AS={5*w_OR_N4*LAMBDA} PS={10*LAMBDA+2*w_OR_N4} AD={5*w_OR_N4*LAMBDA} PD={10*LAMBDA+2*w_OR_N4}

M6      nor       b     gnd   gnd   CMOSN   W={w_OR_N4}   L={2*LAMBDA}
+ AS={5*w_OR_N4*LAMBDA} PS={10*LAMBDA+2*w_OR_N4} AD={5*w_OR_N4*LAMBDA} PD={10*LAMBDA+2*w_OR_N4}

M7      nor       c     gnd   gnd   CMOSN   W={w_OR_N4}   L={2*LAMBDA}
+ AS={5*w_OR_N4*LAMBDA} PS={10*LAMBDA+2*w_OR_N4} AD={5*w_OR_N4*LAMBDA} PD={10*LAMBDA+2*w_OR_N4}

M8      nor       d     gnd   gnd   CMOSN   W={w_OR_N4}   L={2*LAMBDA}
+ AS={5*w_OR_N4*LAMBDA} PS={10*LAMBDA+2*w_OR_N4} AD={5*w_OR_N4*LAMBDA} PD={10*LAMBDA+2*w_OR_N4}

// Inverter
M9      y       nor       vdd     vdd  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

M10      y       nor       gnd     gnd  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
.ends or4_subckt

.subckt and3_subckt a b c y vdd gnd
.param w_AND_P3 = {2*W}
.param w_AND_N3 = {3*W}
//NAND
M1      nand       a       vdd    vdd  CMOSP   W={w_AND_P3}   L={2*LAMBDA}
+ AS={5*w_AND_P3*LAMBDA} PS={10*LAMBDA+2*w_AND_P3} AD={5*w_AND_P3*LAMBDA} PD={10*LAMBDA+2*w_AND_P3}

M2      nand       b       vdd    vdd  CMOSP   W={w_AND_P3}   L={2*LAMBDA}
+ AS={5*w_AND_P3*LAMBDA} PS={10*LAMBDA+2*w_AND_P3} AD={5*w_AND_P3*LAMBDA} PD={10*LAMBDA+2*w_AND_P3}

M3      nand       c       vdd    vdd  CMOSP   W={w_AND_P3}   L={2*LAMBDA}
+ AS={5*w_AND_P3*LAMBDA} PS={10*LAMBDA+2*w_AND_P3} AD={5*w_AND_P3*LAMBDA} PD={10*LAMBDA+2*w_AND_P3}

M4      nand       a       J1     J1   CMOSN   W={w_AND_N3}   L={2*LAMBDA}
+ AS={5*w_AND_N3*LAMBDA} PS={10*LAMBDA+2*w_AND_N3} AD={5*w_AND_N3*LAMBDA} PD={10*LAMBDA+2*w_AND_N3}

M5      J1         b       J2     J2   CMOSN   W={w_AND_N3}   L={2*LAMBDA}
+ AS={5*w_AND_N3*LAMBDA} PS={10*LAMBDA+2*w_AND_N3} AD={5*w_AND_N3*LAMBDA} PD={10*LAMBDA+2*w_AND_N3}

M6      J2         c      gnd    gnd   CMOSN   W={w_AND_N3}   L={2*LAMBDA}
+ AS={5*w_AND_N3*LAMBDA} PS={10*LAMBDA+2*w_AND_N3} AD={5*w_AND_N3*LAMBDA} PD={10*LAMBDA+2*w_AND_N3}

//Inverter
M7      y       nand       vdd     vdd  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

M8      y       nand       gnd     gnd  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
.ends and3_subckt

.subckt and4_subckt a b c d y vdd gnd
.param w_AND_P4 = {2*W}
.param w_AND_N4 = {4*W}
//NAND
M1      nand       a       vdd    vdd  CMOSP   W={w_AND_P4}   L={2*LAMBDA}
+ AS={5*w_AND_P4*LAMBDA} PS={10*LAMBDA+2*w_AND_P4} AD={5*w_AND_P4*LAMBDA} PD={10*LAMBDA+2*w_AND_P4}

M2      nand       b       vdd    vdd  CMOSP   W={w_AND_P4}   L={2*LAMBDA}
+ AS={5*w_AND_P4*LAMBDA} PS={10*LAMBDA+2*w_AND_P4} AD={5*w_AND_P4*LAMBDA} PD={10*LAMBDA+2*w_AND_P4}

M3      nand       c       vdd    vdd  CMOSP   W={w_AND_P4}   L={2*LAMBDA}
+ AS={5*w_AND_N4*LAMBDA} PS={10*LAMBDA+2*w_AND_N4} AD={5*w_AND_N4*LAMBDA} PD={10*LAMBDA+2*w_AND_N4}

M8      J3         d      gnd    gnd   CMOSN   W={w_AND_N4}   L={2*LAMBDA}
+ AS={5*w_AND_N4*LAMBDA} PS={10*LAMBDA+2*w_AND_N4} AD={5*w_AND_N4*LAMBDA} PD={10*LAMBDA+2*w_AND_N4}

//Inverter
M9      y       nand       vdd     vdd  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

M10     y       nand       gnd     gnd  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
.ends and4_subckt




// Carry Calculation
    // Cout1
    // Cout2
        x9  P2 G1 T2_1 vdd gnd and_subckt
        x10 G2 T2_1 Cout2 vdd gnd or_subckt
    // Cout3
        x11 P3 G2 T3_1 vdd gnd and_subckt
        x12 P3 P2 G1 T3_2 vdd gnd and3_subckt
        x13 G3 T3_1 T3_2 Cout3 vdd gnd or3_subckt
    // Cout4
        x14 P4 G3 T4_1 vdd gnd and_subckt
        x15 P4 P3 G2 T4_2 vdd gnd and3_subckt
        x16 P4 P3 P2 G1 T4_3 vdd gnd and4_subckt
        x17 G4 T4_1 T4_2 T4_3 Cout4 vdd gnd or4_subckt



.measure tran rise
+TRIG v(P4) VAL = 0.9V RISE = 1 TARG v(Cout4) VAL = 0.9V RISE = 1
.measure tran FALL
+TRIG v(G4) VAL = 0.9V FALL = 1 TARG v(Cout4) VAL = 0.9V FALL = 1
.measure tran propDelay param='(rise+fall)/2' goal = 0


.tran 1n 200n
.control
set hcopypscolor = 1
set color0=white
set color1=black

run
plot v(G1) v(Cout2)+2  v(Cout3)+4  v(Cout4)+6
set curplottitle= "Aravind Narayanan-2019102014"
plot v(G1) v(G2)+2  v(G3)+4  v(G4)+6
set curplottitle= "Aravind Narayanan-2019102014"
plot v(P1) v(P2)+2  v(P3)+4  v(P4)+6
set curplottitle= "Aravind Narayanan-2019102014"
.endc