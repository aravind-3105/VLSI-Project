* SPICE3 file created from Updated_XOR_WITH.ext - technology: scmos

.option scale=0.09u

M1000 B_bar B 2INV_1/a_6_87# 2INV_1/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1001 B_bar B gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=160 ps=92
M1002 A_bar A vdd 2INV_0/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=340 ps=142
M1003 A_bar A gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1004 vdd A_bar a_56_27# w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=400 ps=180
M1005 a_71_27# B_bar vdd w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1006 out A a_71_27# w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1007 a_56_27# B out w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1008 a_63_n51# A_bar out Gnd nfet w=10 l=2
+  ad=60 pd=32 as=100 ps=60
M1009 gnd B_bar a_63_n51# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1010 a_79_n51# A gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1011 out B a_79_n51# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
C0 a_56_27# out 1.1fF
C1 out gnd! 1.0fF
C2 w_50_21# gnd! 3.0fF
C3 vdd gnd! 3.0fF
C4 gnd gnd! 2.2fF
