magic
tech scmos
timestamp 1619504458
<< nwell >>
rect -16 11 8 43
<< ntransistor >>
rect -5 -7 -3 3
<< ptransistor >>
rect -5 17 -3 37
<< ndiffusion >>
rect -6 -7 -5 3
rect -3 -7 -2 3
<< pdiffusion >>
rect -6 17 -5 37
rect -3 17 -2 37
<< ndcontact >>
rect -10 -7 -6 3
rect -2 -7 2 3
<< pdcontact >>
rect -10 17 -6 37
rect -2 17 2 37
<< polysilicon >>
rect -5 37 -3 40
rect -5 3 -3 17
rect -5 -10 -3 -7
<< polycontact >>
rect -9 6 -5 10
<< metal1 >>
rect -16 42 8 46
rect -10 37 -6 42
rect -2 10 2 17
rect -16 6 -9 10
rect -2 6 8 10
rect -2 3 2 6
rect -10 -11 -6 -7
rect -16 -15 8 -11
<< end >>
