* SPICE3 file created from 4NOR.ext - technology: scmos
.option scale=0.09u
.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.global gnd vdd

Vdd	vdd	gnd	'SUPPLY'
vdA     A     0 pulse 1.8 0 0ns  100ps  100ps 5ns  30ns
vdB     B     0 pulse 1.8 0 30ns 100ps  100ps 10ns  30ns
vdC     C     0 pulse 1.8 0 30ns 100ps  100ps 20ns  40ns
vd4     D     0 pulse 1.8 0 2ns  100ps  100ps 30ns  50ns

M1000 a_13_6# D vdd w_0_0# CMOSP w=80 l=2
+  ad=480 pd=172 as=400 ps=170
M1001 a_21_6# C a_13_6# w_0_0# CMOSP w=80 l=2
+  ad=480 pd=172 as=0 ps=0
M1002 a_29_6# B a_21_6# w_0_0# CMOSP w=80 l=2
+  ad=480 pd=172 as=0 ps=0
M1003 out A a_29_6# w_0_0# CMOSP w=80 l=2
+  ad=560 pd=174 as=0 ps=0
M1004 out D gnd gnd CMOSN w=10 l=2
+  ad=120 pd=64 as=180 ps=96
M1005 gnd C out gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 out B gnd gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 gnd A out gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
C0 w_0_0# gnd 4.9fF



.tran 1n 60n
.control
set hcopypscolor = 1
set color0=white
set color1=black

run
plot v(A) v(B)+2 v(C)+4 v(D)+8 v(out)+10
set curplottitle= "Aravind Narayanan-2019102014"
.endc