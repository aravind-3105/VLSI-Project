magic
tech scmos
timestamp 1619551394
<< metal1 >>
rect -34 -95 -29 140
rect -23 35 -18 158
rect -10 42 -5 122
rect -10 38 3 42
rect 60 38 82 42
rect -23 31 3 35
rect 1 0 3 4
rect 77 -7 82 38
rect -9 -12 82 -7
rect -9 -88 -4 -12
rect -9 -92 6 -88
rect -34 -99 4 -95
rect 62 -108 79 -104
rect 3 -129 6 -125
rect 73 -145 79 -108
rect 216 -133 221 172
rect 231 120 236 184
rect 232 36 236 120
rect 243 43 247 141
rect 348 47 352 183
rect 359 55 363 158
rect 368 62 372 121
rect 368 58 382 62
rect 445 59 467 63
rect 359 50 381 55
rect 348 43 382 47
rect 243 39 251 43
rect 309 39 331 43
rect 232 32 257 36
rect 326 -126 331 39
rect 374 1 386 5
rect 462 -7 467 59
rect 361 -12 467 -7
rect 361 -119 367 -12
rect 361 -123 380 -119
rect 326 -130 386 -126
rect 216 -137 389 -133
rect 447 -144 483 -140
rect 72 -201 79 -145
rect 378 -165 389 -161
rect 477 -201 483 -144
rect 574 -155 580 208
rect 742 202 747 203
rect 870 202 875 203
rect 605 36 611 196
rect 621 43 626 173
rect 742 47 747 196
rect 754 55 759 183
rect 766 62 771 141
rect 766 58 782 62
rect 843 59 857 63
rect 754 51 782 55
rect 742 43 786 47
rect 621 39 639 43
rect 694 39 719 43
rect 605 32 642 36
rect 713 -148 719 39
rect 778 1 786 5
rect 853 -141 857 59
rect 870 57 875 196
rect 884 64 889 183
rect 897 71 902 157
rect 908 128 912 132
rect 908 78 912 122
rect 908 74 923 78
rect 995 74 1014 78
rect 897 67 926 71
rect 884 60 934 64
rect 870 53 936 57
rect 916 2 929 6
rect 902 -6 907 -5
rect 1009 -6 1014 74
rect 902 -11 1014 -6
rect 902 -134 907 -11
rect 902 -138 914 -134
rect 853 -145 922 -141
rect 713 -152 921 -148
rect 574 -159 916 -155
rect 990 -166 1047 -162
rect 915 -187 926 -182
rect 1043 -234 1047 -166
<< m2contact >>
rect 574 208 580 215
rect 231 184 236 190
rect 215 172 222 178
rect -23 158 -18 165
rect -34 140 -28 147
rect -10 122 -3 130
rect -1 73 7 82
rect 57 74 63 79
rect -4 0 1 5
rect 57 -72 63 -67
rect -2 -129 3 -123
rect 57 -134 63 -125
rect 348 183 353 189
rect 243 141 249 148
rect 250 76 257 83
rect 307 75 314 80
rect 359 158 364 165
rect 368 121 374 129
rect 376 95 383 100
rect 440 95 448 101
rect 308 16 314 22
rect 368 1 374 7
rect 443 -108 451 -102
rect 373 -165 378 -159
rect 442 -168 449 -161
rect 605 196 612 202
rect 741 196 748 202
rect 869 196 876 202
rect 621 173 628 179
rect 633 76 640 82
rect 691 75 697 81
rect 754 183 760 189
rect 766 141 773 147
rect 775 95 781 101
rect 839 95 845 101
rect 688 17 696 23
rect 839 37 846 43
rect 771 0 778 6
rect 884 183 890 190
rect 897 157 903 165
rect 908 122 914 128
rect 916 110 922 116
rect 990 110 997 116
rect 910 1 916 7
rect 988 -129 995 -124
rect 907 -187 915 -180
<< metal2 >>
rect -190 -142 -181 227
rect -109 210 574 215
rect -110 197 605 202
rect 612 197 741 202
rect 748 197 869 202
rect -110 184 231 188
rect 236 184 348 188
rect -110 183 348 184
rect 353 183 754 188
rect 760 183 884 188
rect 890 183 891 188
rect -109 173 215 178
rect 222 173 621 178
rect -108 158 -23 164
rect -18 158 359 164
rect 364 158 897 164
rect -109 141 -34 146
rect -28 141 243 146
rect 249 141 766 146
rect -109 122 -10 127
rect -3 122 368 127
rect 374 122 908 127
rect 374 121 913 122
rect 841 111 916 115
rect 635 101 641 102
rect 841 101 846 111
rect 997 110 1028 115
rect 308 95 376 100
rect 482 100 641 101
rect 448 95 641 100
rect -105 75 -1 81
rect 92 79 250 81
rect 63 76 250 79
rect 308 80 313 95
rect 63 75 254 76
rect -17 0 -4 4
rect -17 -124 -13 0
rect 92 -68 96 75
rect 63 -72 96 -68
rect 309 6 313 16
rect 309 1 368 6
rect -110 -129 -2 -124
rect -110 -130 3 -129
rect 309 -128 313 1
rect 482 -103 488 95
rect 635 82 641 95
rect 640 80 641 82
rect 692 95 775 100
rect 845 96 846 101
rect 692 94 779 95
rect 692 81 698 94
rect 697 76 698 81
rect 910 43 915 44
rect 846 38 915 43
rect 696 17 777 22
rect 689 16 777 17
rect 451 -108 488 -103
rect 63 -134 314 -128
rect 309 -159 313 -134
rect 309 -163 373 -159
rect 691 -162 696 16
rect 771 6 777 16
rect 910 7 915 38
rect 1023 -74 1028 110
rect 988 -79 1028 -74
rect 988 -124 992 -79
rect 449 -168 697 -162
rect 691 -180 696 -168
rect 691 -186 907 -180
use and2  and2_0
timestamp 1619509263
transform 1 0 46 0 1 -12
box -46 12 16 90
use and2  and2_1
timestamp 1619509263
transform 1 0 296 0 1 -11
box -46 12 16 90
use and3  and3_0
timestamp 1619507409
transform 1 0 422 0 1 38
box -46 -37 24 61
use and2  and2_2
timestamp 1619509263
transform 1 0 679 0 1 -11
box -46 12 16 90
use and3  and3_1
timestamp 1619507409
transform 1 0 821 0 1 38
box -46 -37 24 61
use and4  and4_0
timestamp 1619509145
transform 1 0 971 0 1 53
box -54 -51 24 61
use or2  or2_0
timestamp 1619513079
transform 1 0 38 0 1 -129
box -38 0 24 97
use or3  or3_0
timestamp 1619513799
transform 1 0 424 0 1 -165
box -46 0 24 122
use or4  or4_0
timestamp 1619514549
transform 1 0 968 0 1 -187
box -56 0 24 149
<< labels >>
rlabel metal2 -94 -127 -94 -127 1 gnd
rlabel metal2 -93 78 -93 78 1 vdd
rlabel metal2 -93 125 -93 125 1 g1
rlabel metal2 -95 143 -95 143 1 g2
rlabel metal2 -95 160 -95 160 1 p2
rlabel metal2 -96 176 -96 176 1 g3
rlabel metal2 -96 186 -96 186 1 p3
rlabel metal2 -98 200 -98 200 1 p4
rlabel metal2 -97 213 -97 213 1 g4
rlabel metal1 76 -177 76 -177 1 c2
rlabel metal1 480 -188 480 -188 1 c3
rlabel metal1 1045 -208 1045 -208 7 c4
rlabel metal2 -186 214 -186 214 3 g1
rlabel metal2 -186 -126 -186 -126 3 c1
<< end >>
