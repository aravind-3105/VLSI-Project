magic
tech scmos
timestamp 1619560144
<< nwell >>
rect 50 21 98 77
<< ntransistor >>
rect 61 -51 63 -41
rect 69 -51 71 -41
rect 77 -51 79 -41
rect 85 -51 87 -41
<< ptransistor >>
rect 61 27 63 67
rect 69 27 71 67
rect 77 27 79 67
rect 85 27 87 67
<< ndiffusion >>
rect 60 -51 61 -41
rect 63 -51 69 -41
rect 71 -51 72 -41
rect 76 -51 77 -41
rect 79 -51 85 -41
rect 87 -51 88 -41
<< pdiffusion >>
rect 60 27 61 67
rect 63 27 64 67
rect 68 27 69 67
rect 71 27 72 67
rect 76 27 77 67
rect 79 27 80 67
rect 84 27 85 67
rect 87 27 88 67
<< ndcontact >>
rect 56 -51 60 -41
rect 72 -51 76 -41
rect 88 -51 92 -41
<< pdcontact >>
rect 6 42 10 62
rect 56 27 60 67
rect 64 27 68 67
rect 72 27 76 67
rect 80 27 84 67
rect 88 27 92 67
<< polysilicon >>
rect 61 67 63 70
rect 69 67 71 70
rect 77 67 79 70
rect 85 67 87 70
rect 61 3 63 27
rect 61 -11 63 -1
rect 51 -13 63 -11
rect 51 -57 53 -13
rect 69 -20 71 27
rect 77 18 79 27
rect 61 -22 71 -20
rect 61 -26 63 -22
rect 61 -41 63 -30
rect 69 -41 71 -38
rect 77 -41 79 14
rect 85 11 87 27
rect 85 -41 87 7
rect 61 -54 63 -51
rect 69 -57 71 -51
rect 77 -54 79 -51
rect 85 -54 87 -51
rect 51 -59 71 -57
<< polycontact >>
rect 59 -1 63 3
rect 75 14 79 18
rect 59 -30 63 -26
rect 83 7 87 11
<< metal1 >>
rect 20 73 68 77
rect 20 71 24 73
rect -1 66 24 71
rect 64 67 68 73
rect 80 73 99 77
rect 80 67 84 73
rect -20 29 6 33
rect -8 -3 -4 29
rect 21 23 34 27
rect 56 24 60 27
rect 88 24 92 27
rect 56 21 92 24
rect 43 14 75 18
rect 43 -3 47 14
rect 95 11 99 73
rect -8 -7 47 -3
rect 50 7 83 11
rect 90 7 99 11
rect 50 -10 53 7
rect -15 -14 53 -10
rect 56 -1 59 3
rect -15 -59 -11 -14
rect 56 -18 60 -1
rect -1 -26 24 -21
rect 90 -9 94 7
rect 90 -13 103 -9
rect 41 -30 59 -26
rect -20 -63 5 -59
rect 41 -65 45 -30
rect 90 -33 94 -13
rect 72 -36 94 -33
rect 72 -41 76 -36
rect 18 -69 45 -65
rect 56 -87 60 -51
rect -15 -92 24 -87
rect 29 -88 60 -87
rect 88 -88 92 -51
rect 29 -92 92 -88
<< m2contact >>
rect -6 66 -1 71
rect 34 23 39 28
rect 22 0 27 5
rect -6 -26 -1 -21
rect 55 -23 60 -18
rect 24 -92 29 -87
<< metal2 >>
rect -6 -21 -2 66
rect 23 -16 27 0
rect 23 -20 29 -16
rect 25 -87 29 -20
rect 35 -18 39 23
rect 35 -23 55 -18
use 2INV  2INV_0
timestamp 1619542334
transform 1 0 0 0 1 -45
box 0 45 24 116
use 2INV  2INV_1
timestamp 1619542334
transform 1 0 0 0 1 -137
box 0 45 24 116
<< end >>
