magic
tech scmos
timestamp 1619455295
<< nwell >>
rect 0 0 52 32
<< ntransistor >>
rect 11 -78 13 -38
rect 19 -78 21 -38
rect 27 -78 29 -38
rect 35 -78 37 -38
<< ptransistor >>
rect 11 6 13 26
rect 19 6 21 26
rect 27 6 29 26
rect 35 6 37 26
<< ndiffusion >>
rect 10 -78 11 -38
rect 13 -78 19 -38
rect 21 -78 27 -38
rect 29 -78 35 -38
rect 37 -78 40 -38
<< pdiffusion >>
rect 10 6 11 26
rect 13 6 14 26
rect 18 6 19 26
rect 21 6 22 26
rect 26 6 27 26
rect 29 6 30 26
rect 34 6 35 26
rect 37 6 38 26
<< ndcontact >>
rect 6 -78 10 -38
rect 40 -78 44 -38
<< pdcontact >>
rect 6 6 10 26
rect 14 6 18 26
rect 22 6 26 26
rect 30 6 34 26
rect 38 6 42 26
<< polysilicon >>
rect 11 26 13 29
rect 19 26 21 29
rect 27 26 29 29
rect 35 26 37 29
rect 11 -31 13 6
rect 19 -24 21 6
rect 27 -17 29 6
rect 35 -10 37 6
rect 11 -38 13 -35
rect 19 -38 21 -28
rect 27 -38 29 -21
rect 35 -38 37 -14
rect 11 -82 13 -78
rect 19 -82 21 -78
rect 27 -82 29 -78
rect 35 -82 37 -78
<< polycontact >>
rect 33 -14 37 -10
rect 25 -21 29 -17
rect 17 -28 21 -24
rect 9 -35 13 -31
<< metal1 >>
rect 0 30 52 33
rect 6 26 10 30
rect 22 26 26 30
rect 38 26 42 30
rect 14 -3 18 6
rect 30 -3 34 6
rect 14 -7 52 -3
rect 0 -14 33 -10
rect 0 -21 25 -17
rect 0 -28 17 -24
rect 0 -35 9 -31
rect 40 -38 44 -7
rect 6 -83 10 -78
rect 0 -86 52 -83
<< labels >>
rlabel metal1 2 -12 2 -12 3 A
rlabel metal1 2 -19 2 -19 3 B
rlabel metal1 2 -26 2 -26 3 C
rlabel metal1 2 -33 2 -33 3 D
rlabel metal1 48 -5 48 -5 7 out
rlabel metal1 25 -85 25 -85 1 gnd
rlabel metal1 24 32 24 32 5 vdd
<< end >>
