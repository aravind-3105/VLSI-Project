* SPICE3 file created from 2AND_WI.ext - technology: scmos

.option scale=0.01u

M1000 out out_bar 2INV_0/a_6_87# 2INV_0/w_0_81# pfet w=180 l=18
+  ad=8100 pd=450 as=8100 ps=450
M1001 out out_bar gnd Gnd nfet w=90 l=18
+  ad=4050 pd=270 as=12150 ps=720
M1002 out_bar A vdd 2NAND_WO_0/w_0_0# pfet w=180 l=18
+  ad=9720 pd=468 as=16200 ps=900
M1003 vdd B out_bar 2NAND_WO_0/w_0_0# pfet w=180 l=18
+  ad=0 pd=0 as=0 ps=0
M1004 2NAND_WO_0/a_13_n43# A gnd Gnd nfet w=180 l=18
+  ad=9720 pd=468 as=0 ps=0
M1005 out_bar B 2NAND_WO_0/a_13_n43# Gnd nfet w=180 l=18
+  ad=11340 pd=486 as=0 ps=0
C0 2NAND_WO_0/w_0_0# gnd! 1.2fF
