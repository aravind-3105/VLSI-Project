* SPICE3 file created from FullBlock_WI_Updated.ext - technology: scmos

.option scale=0.09u

M1000 SUM_WO_0/XOR_WO_3/a_59_n30# c3 SUM_WO_0/XOR_WO_3/2INV_1/a_6_87# SUM_WO_0/XOR_WO_3/2INV_1/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1001 SUM_WO_0/XOR_WO_3/a_59_n30# c3 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=3840 ps=2148
M1002 SUM_WO_0/XOR_WO_3/a_51_n59# p4 vdd SUM_WO_0/XOR_WO_3/2INV_0/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=5780 ps=2582
M1003 SUM_WO_0/XOR_WO_3/a_51_n59# p4 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1004 vdd SUM_WO_0/XOR_WO_3/a_51_n59# SUM_WO_0/XOR_WO_3/a_56_27# SUM_WO_0/XOR_WO_3/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=400 ps=180
M1005 SUM_WO_0/XOR_WO_3/a_71_27# SUM_WO_0/XOR_WO_3/a_59_n30# vdd SUM_WO_0/XOR_WO_3/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1006 s4 p4 SUM_WO_0/XOR_WO_3/a_71_27# SUM_WO_0/XOR_WO_3/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1007 SUM_WO_0/XOR_WO_3/a_56_27# c3 s4 SUM_WO_0/XOR_WO_3/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1008 SUM_WO_0/XOR_WO_3/a_63_n51# SUM_WO_0/XOR_WO_3/a_59_n30# gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1009 s4 SUM_WO_0/XOR_WO_3/a_51_n59# SUM_WO_0/XOR_WO_3/a_63_n51# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1010 SUM_WO_0/XOR_WO_3/a_79_n51# p4 s4 Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1011 gnd c3 SUM_WO_0/XOR_WO_3/a_79_n51# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1012 SUM_WO_0/XOR_WO_2/a_59_n30# c2 SUM_WO_0/XOR_WO_2/2INV_1/a_6_87# SUM_WO_0/XOR_WO_2/2INV_1/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1013 SUM_WO_0/XOR_WO_2/a_59_n30# c2 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1014 SUM_WO_0/XOR_WO_2/a_51_n59# p3 vdd SUM_WO_0/XOR_WO_2/2INV_0/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1015 SUM_WO_0/XOR_WO_2/a_51_n59# p3 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1016 vdd SUM_WO_0/XOR_WO_2/a_51_n59# SUM_WO_0/XOR_WO_2/a_56_27# SUM_WO_0/XOR_WO_2/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=400 ps=180
M1017 SUM_WO_0/XOR_WO_2/a_71_27# SUM_WO_0/XOR_WO_2/a_59_n30# vdd SUM_WO_0/XOR_WO_2/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1018 s3 p3 SUM_WO_0/XOR_WO_2/a_71_27# SUM_WO_0/XOR_WO_2/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1019 SUM_WO_0/XOR_WO_2/a_56_27# c2 s3 SUM_WO_0/XOR_WO_2/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1020 SUM_WO_0/XOR_WO_2/a_63_n51# SUM_WO_0/XOR_WO_2/a_59_n30# gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1021 s3 SUM_WO_0/XOR_WO_2/a_51_n59# SUM_WO_0/XOR_WO_2/a_63_n51# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1022 SUM_WO_0/XOR_WO_2/a_79_n51# p3 s3 Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1023 gnd c2 SUM_WO_0/XOR_WO_2/a_79_n51# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1024 SUM_WO_0/XOR_WO_1/a_59_n30# g1 SUM_WO_0/XOR_WO_1/2INV_1/a_6_87# SUM_WO_0/XOR_WO_1/2INV_1/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1025 SUM_WO_0/XOR_WO_1/a_59_n30# g1 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1026 SUM_WO_0/XOR_WO_1/a_51_n59# p2 vdd SUM_WO_0/XOR_WO_1/2INV_0/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1027 SUM_WO_0/XOR_WO_1/a_51_n59# p2 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1028 vdd SUM_WO_0/XOR_WO_1/a_51_n59# SUM_WO_0/XOR_WO_1/a_56_27# SUM_WO_0/XOR_WO_1/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=400 ps=180
M1029 SUM_WO_0/XOR_WO_1/a_71_27# SUM_WO_0/XOR_WO_1/a_59_n30# vdd SUM_WO_0/XOR_WO_1/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1030 s2 p2 SUM_WO_0/XOR_WO_1/a_71_27# SUM_WO_0/XOR_WO_1/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1031 SUM_WO_0/XOR_WO_1/a_56_27# g1 s2 SUM_WO_0/XOR_WO_1/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1032 SUM_WO_0/XOR_WO_1/a_63_n51# SUM_WO_0/XOR_WO_1/a_59_n30# gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1033 s2 SUM_WO_0/XOR_WO_1/a_51_n59# SUM_WO_0/XOR_WO_1/a_63_n51# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1034 SUM_WO_0/XOR_WO_1/a_79_n51# p2 s2 Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1035 gnd g1 SUM_WO_0/XOR_WO_1/a_79_n51# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1036 SUM_WO_0/XOR_WO_0/a_59_n30# gnd SUM_WO_0/XOR_WO_0/2INV_1/a_6_87# SUM_WO_0/XOR_WO_0/2INV_1/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1037 SUM_WO_0/XOR_WO_0/a_59_n30# gnd gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1038 SUM_WO_0/XOR_WO_0/a_51_n59# p1 vdd SUM_WO_0/XOR_WO_0/2INV_0/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1039 SUM_WO_0/XOR_WO_0/a_51_n59# p1 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1040 vdd SUM_WO_0/XOR_WO_0/a_51_n59# SUM_WO_0/XOR_WO_0/a_56_27# SUM_WO_0/XOR_WO_0/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=400 ps=180
M1041 SUM_WO_0/XOR_WO_0/a_71_27# SUM_WO_0/XOR_WO_0/a_59_n30# vdd SUM_WO_0/XOR_WO_0/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1042 s1 p1 SUM_WO_0/XOR_WO_0/a_71_27# SUM_WO_0/XOR_WO_0/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1043 SUM_WO_0/XOR_WO_0/a_56_27# gnd s1 SUM_WO_0/XOR_WO_0/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1044 SUM_WO_0/XOR_WO_0/a_63_n51# SUM_WO_0/XOR_WO_0/a_59_n30# gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1045 s1 SUM_WO_0/XOR_WO_0/a_51_n59# SUM_WO_0/XOR_WO_0/a_63_n51# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1046 SUM_WO_0/XOR_WO_0/a_79_n51# p1 s1 Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1047 gnd gnd SUM_WO_0/XOR_WO_0/a_79_n51# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1048 c4 Carry_WO_0/m1_409_n151# Carry_WO_0/2INV_8/a_6_87# Carry_WO_0/2INV_8/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1049 c4 Carry_WO_0/m1_409_n151# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1050 Carry_WO_0/4NOR_WO_0/a_13_6# Carry_WO_0/m1_395_n85# vdd Carry_WO_0/4NOR_WO_0/w_0_0# pfet w=80 l=2
+  ad=480 pd=172 as=0 ps=0
M1051 Carry_WO_0/4NOR_WO_0/a_21_6# Carry_WO_0/m1_402_n83# Carry_WO_0/4NOR_WO_0/a_13_6# Carry_WO_0/4NOR_WO_0/w_0_0# pfet w=80 l=2
+  ad=480 pd=172 as=0 ps=0
M1052 Carry_WO_0/4NOR_WO_0/a_29_6# Carry_WO_0/m1_409_n82# Carry_WO_0/4NOR_WO_0/a_21_6# Carry_WO_0/4NOR_WO_0/w_0_0# pfet w=80 l=2
+  ad=480 pd=172 as=0 ps=0
M1053 Carry_WO_0/m1_409_n151# g4 Carry_WO_0/4NOR_WO_0/a_29_6# Carry_WO_0/4NOR_WO_0/w_0_0# pfet w=80 l=2
+  ad=560 pd=174 as=0 ps=0
M1054 Carry_WO_0/m1_409_n151# Carry_WO_0/m1_395_n85# gnd Gnd nfet w=10 l=2
+  ad=120 pd=64 as=0 ps=0
M1055 gnd Carry_WO_0/m1_402_n83# Carry_WO_0/m1_409_n151# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1056 Carry_WO_0/m1_409_n151# Carry_WO_0/m1_409_n82# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1057 gnd g4 Carry_WO_0/m1_409_n151# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1058 Carry_WO_0/m1_409_n82# Carry_WO_0/m1_683_20# Carry_WO_0/2INV_7/a_6_87# Carry_WO_0/2INV_7/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1059 Carry_WO_0/m1_409_n82# Carry_WO_0/m1_683_20# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1060 Carry_WO_0/m1_683_20# p4 vdd Carry_WO_0/4NAND_WO_0/w_0_0# pfet w=20 l=2
+  ad=240 pd=104 as=0 ps=0
M1061 vdd p3 Carry_WO_0/m1_683_20# Carry_WO_0/4NAND_WO_0/w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1062 Carry_WO_0/m1_683_20# p2 vdd Carry_WO_0/4NAND_WO_0/w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1063 vdd g1 Carry_WO_0/m1_683_20# Carry_WO_0/4NAND_WO_0/w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1064 Carry_WO_0/4NAND_WO_0/a_13_n78# p4 gnd Gnd nfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1065 Carry_WO_0/4NAND_WO_0/a_21_n78# p3 Carry_WO_0/4NAND_WO_0/a_13_n78# Gnd nfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1066 Carry_WO_0/4NAND_WO_0/a_29_n78# p2 Carry_WO_0/4NAND_WO_0/a_21_n78# Gnd nfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1067 Carry_WO_0/m1_683_20# g1 Carry_WO_0/4NAND_WO_0/a_29_n78# Gnd nfet w=40 l=2
+  ad=280 pd=94 as=0 ps=0
M1068 Carry_WO_0/3NOR_WO_0/a_14_3# Carry_WO_0/m1_174_23# vdd Carry_WO_0/3NOR_WO_0/w_1_n3# pfet w=60 l=2
+  ad=360 pd=132 as=0 ps=0
M1069 Carry_WO_0/3NOR_WO_0/a_22_3# g3 Carry_WO_0/3NOR_WO_0/a_14_3# Carry_WO_0/3NOR_WO_0/w_1_n3# pfet w=60 l=2
+  ad=360 pd=132 as=0 ps=0
M1070 Carry_WO_0/m1_194_n80# Carry_WO_0/m1_226_n94# Carry_WO_0/3NOR_WO_0/a_22_3# Carry_WO_0/3NOR_WO_0/w_1_n3# pfet w=60 l=2
+  ad=420 pd=134 as=0 ps=0
M1071 Carry_WO_0/m1_194_n80# Carry_WO_0/m1_174_23# gnd Gnd nfet w=10 l=2
+  ad=130 pd=66 as=0 ps=0
M1072 gnd g3 Carry_WO_0/m1_194_n80# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1073 Carry_WO_0/m1_194_n80# Carry_WO_0/m1_226_n94# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1074 c3 Carry_WO_0/m1_194_n80# Carry_WO_0/2INV_3/a_6_87# Carry_WO_0/2INV_3/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1075 c3 Carry_WO_0/m1_194_n80# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1076 Carry_WO_0/m1_402_n83# Carry_WO_0/m1_526_53# Carry_WO_0/2INV_6/a_6_87# Carry_WO_0/2INV_6/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1077 Carry_WO_0/m1_402_n83# Carry_WO_0/m1_526_53# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1078 Carry_WO_0/m1_526_53# p4 vdd Carry_WO_0/3NAND_WO_1/w_0_0# pfet w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M1079 vdd p3 Carry_WO_0/m1_526_53# Carry_WO_0/3NAND_WO_1/w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1080 Carry_WO_0/m1_526_53# g2 vdd Carry_WO_0/3NAND_WO_1/w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1081 Carry_WO_0/3NAND_WO_1/a_13_n61# p4 gnd Gnd nfet w=30 l=2
+  ad=180 pd=72 as=0 ps=0
M1082 Carry_WO_0/3NAND_WO_1/a_21_n61# p3 Carry_WO_0/3NAND_WO_1/a_13_n61# Gnd nfet w=30 l=2
+  ad=180 pd=72 as=0 ps=0
M1083 Carry_WO_0/m1_526_53# g2 Carry_WO_0/3NAND_WO_1/a_21_n61# Gnd nfet w=30 l=2
+  ad=210 pd=74 as=0 ps=0
M1084 Carry_WO_0/m1_395_n85# Carry_WO_0/m1_398_36# Carry_WO_0/2INV_5/a_6_87# Carry_WO_0/2INV_5/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1085 Carry_WO_0/m1_395_n85# Carry_WO_0/m1_398_36# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1086 Carry_WO_0/m1_398_36# p4 vdd Carry_WO_0/2NAND_WO_2/w_0_0# pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1087 vdd g3 Carry_WO_0/m1_398_36# Carry_WO_0/2NAND_WO_2/w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1088 Carry_WO_0/2NAND_WO_2/a_13_n43# p4 gnd Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1089 Carry_WO_0/m1_398_36# g3 Carry_WO_0/2NAND_WO_2/a_13_n43# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1090 Carry_WO_0/m1_226_n94# Carry_WO_0/m1_252_46# Carry_WO_0/2INV_4/a_6_87# Carry_WO_0/2INV_4/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1091 Carry_WO_0/m1_226_n94# Carry_WO_0/m1_252_46# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1092 Carry_WO_0/m1_252_46# g1 vdd Carry_WO_0/3NAND_WO_0/w_0_0# pfet w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M1093 vdd p2 Carry_WO_0/m1_252_46# Carry_WO_0/3NAND_WO_0/w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1094 Carry_WO_0/m1_252_46# p3 vdd Carry_WO_0/3NAND_WO_0/w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1095 Carry_WO_0/3NAND_WO_0/a_13_n61# g1 gnd Gnd nfet w=30 l=2
+  ad=180 pd=72 as=0 ps=0
M1096 Carry_WO_0/3NAND_WO_0/a_21_n61# p2 Carry_WO_0/3NAND_WO_0/a_13_n61# Gnd nfet w=30 l=2
+  ad=180 pd=72 as=0 ps=0
M1097 Carry_WO_0/m1_252_46# p3 Carry_WO_0/3NAND_WO_0/a_21_n61# Gnd nfet w=30 l=2
+  ad=210 pd=74 as=0 ps=0
M1098 Carry_WO_0/m1_174_23# Carry_WO_0/m1_145_29# Carry_WO_0/2INV_2/a_6_87# Carry_WO_0/2INV_2/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1099 Carry_WO_0/m1_174_23# Carry_WO_0/m1_145_29# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1100 Carry_WO_0/m1_145_29# p3 vdd Carry_WO_0/2NAND_WO_1/w_0_0# pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1101 vdd g2 Carry_WO_0/m1_145_29# Carry_WO_0/2NAND_WO_1/w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1102 Carry_WO_0/2NAND_WO_1/a_13_n43# p3 gnd Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1103 Carry_WO_0/m1_145_29# g2 Carry_WO_0/2NAND_WO_1/a_13_n43# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1104 Carry_WO_0/2NOR_WO_0/a_13_5# Carry_WO_0/m1_63_n31# vdd Carry_WO_0/w_38_n91# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1105 Carry_WO_0/m1_19_n37# g2 Carry_WO_0/2NOR_WO_0/a_13_5# Carry_WO_0/w_38_n91# pfet w=40 l=2
+  ad=280 pd=94 as=0 ps=0
M1106 Carry_WO_0/m1_19_n37# Carry_WO_0/m1_63_n31# gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1107 gnd g2 Carry_WO_0/m1_19_n37# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1108 c2 Carry_WO_0/m1_19_n37# Carry_WO_0/2INV_1/a_6_87# Carry_WO_0/2INV_1/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1109 c2 Carry_WO_0/m1_19_n37# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1110 Carry_WO_0/m1_63_n31# Carry_WO_0/m1_25_30# Carry_WO_0/2INV_0/a_6_87# Carry_WO_0/2INV_0/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1111 Carry_WO_0/m1_63_n31# Carry_WO_0/m1_25_30# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1112 Carry_WO_0/m1_25_30# g1 vdd Carry_WO_0/w_7_77# pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1113 vdd p2 Carry_WO_0/m1_25_30# Carry_WO_0/w_7_77# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1114 Carry_WO_0/2NAND_WO_0/a_13_n43# g1 gnd Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1115 Carry_WO_0/m1_25_30# p2 Carry_WO_0/2NAND_WO_0/a_13_n43# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1116 g2 g2_bar PropagateGenerate_WO_0/2INV_3/a_6_87# PropagateGenerate_WO_0/2INV_3/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1117 g2 g2_bar gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1118 g1 g1_bar PropagateGenerate_WO_0/2INV_2/a_6_87# PropagateGenerate_WO_0/2INV_2/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1119 g1 g1_bar gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1120 g3 g3_bar PropagateGenerate_WO_0/2INV_1/a_6_87# PropagateGenerate_WO_0/2INV_1/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1121 g3 g3_bar gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1122 g4 g4_bar PropagateGenerate_WO_0/2INV_0/a_6_87# PropagateGenerate_WO_0/2INV_0/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1123 g4 g4_bar gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1124 PropagateGenerate_WO_0/XOR_WO_3/a_59_n30# b4 PropagateGenerate_WO_0/XOR_WO_3/2INV_1/a_6_87# PropagateGenerate_WO_0/XOR_WO_3/2INV_1/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1125 PropagateGenerate_WO_0/XOR_WO_3/a_59_n30# b4 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1126 PropagateGenerate_WO_0/XOR_WO_3/a_51_n59# a4 vdd PropagateGenerate_WO_0/XOR_WO_3/2INV_0/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1127 PropagateGenerate_WO_0/XOR_WO_3/a_51_n59# a4 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1128 vdd PropagateGenerate_WO_0/XOR_WO_3/a_51_n59# PropagateGenerate_WO_0/XOR_WO_3/a_56_27# PropagateGenerate_WO_0/XOR_WO_3/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=400 ps=180
M1129 PropagateGenerate_WO_0/XOR_WO_3/a_71_27# PropagateGenerate_WO_0/XOR_WO_3/a_59_n30# vdd PropagateGenerate_WO_0/XOR_WO_3/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1130 p4 a4 PropagateGenerate_WO_0/XOR_WO_3/a_71_27# PropagateGenerate_WO_0/XOR_WO_3/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1131 PropagateGenerate_WO_0/XOR_WO_3/a_56_27# b4 p4 PropagateGenerate_WO_0/XOR_WO_3/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1132 PropagateGenerate_WO_0/XOR_WO_3/a_63_n51# PropagateGenerate_WO_0/XOR_WO_3/a_59_n30# gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1133 p4 PropagateGenerate_WO_0/XOR_WO_3/a_51_n59# PropagateGenerate_WO_0/XOR_WO_3/a_63_n51# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1134 PropagateGenerate_WO_0/XOR_WO_3/a_79_n51# a4 p4 Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1135 gnd b4 PropagateGenerate_WO_0/XOR_WO_3/a_79_n51# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1136 PropagateGenerate_WO_0/XOR_WO_2/a_59_n30# b3 PropagateGenerate_WO_0/XOR_WO_2/2INV_1/a_6_87# PropagateGenerate_WO_0/XOR_WO_2/2INV_1/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1137 PropagateGenerate_WO_0/XOR_WO_2/a_59_n30# b3 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1138 PropagateGenerate_WO_0/XOR_WO_2/a_51_n59# a3 vdd PropagateGenerate_WO_0/XOR_WO_2/2INV_0/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1139 PropagateGenerate_WO_0/XOR_WO_2/a_51_n59# a3 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1140 vdd PropagateGenerate_WO_0/XOR_WO_2/a_51_n59# PropagateGenerate_WO_0/XOR_WO_2/a_56_27# PropagateGenerate_WO_0/XOR_WO_2/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=400 ps=180
M1141 PropagateGenerate_WO_0/XOR_WO_2/a_71_27# PropagateGenerate_WO_0/XOR_WO_2/a_59_n30# vdd PropagateGenerate_WO_0/XOR_WO_2/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1142 p3 a3 PropagateGenerate_WO_0/XOR_WO_2/a_71_27# PropagateGenerate_WO_0/XOR_WO_2/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1143 PropagateGenerate_WO_0/XOR_WO_2/a_56_27# b3 p3 PropagateGenerate_WO_0/XOR_WO_2/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1144 PropagateGenerate_WO_0/XOR_WO_2/a_63_n51# PropagateGenerate_WO_0/XOR_WO_2/a_59_n30# gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1145 p3 PropagateGenerate_WO_0/XOR_WO_2/a_51_n59# PropagateGenerate_WO_0/XOR_WO_2/a_63_n51# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1146 PropagateGenerate_WO_0/XOR_WO_2/a_79_n51# a3 p3 Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1147 gnd b3 PropagateGenerate_WO_0/XOR_WO_2/a_79_n51# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1148 PropagateGenerate_WO_0/XOR_WO_1/a_59_n30# b2 PropagateGenerate_WO_0/XOR_WO_1/2INV_1/a_6_87# PropagateGenerate_WO_0/XOR_WO_1/2INV_1/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1149 PropagateGenerate_WO_0/XOR_WO_1/a_59_n30# b2 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1150 PropagateGenerate_WO_0/XOR_WO_1/a_51_n59# a2 vdd PropagateGenerate_WO_0/XOR_WO_1/2INV_0/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1151 PropagateGenerate_WO_0/XOR_WO_1/a_51_n59# a2 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1152 vdd PropagateGenerate_WO_0/XOR_WO_1/a_51_n59# PropagateGenerate_WO_0/XOR_WO_1/a_56_27# PropagateGenerate_WO_0/XOR_WO_1/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=400 ps=180
M1153 PropagateGenerate_WO_0/XOR_WO_1/a_71_27# PropagateGenerate_WO_0/XOR_WO_1/a_59_n30# vdd PropagateGenerate_WO_0/XOR_WO_1/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1154 p2 a2 PropagateGenerate_WO_0/XOR_WO_1/a_71_27# PropagateGenerate_WO_0/XOR_WO_1/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1155 PropagateGenerate_WO_0/XOR_WO_1/a_56_27# b2 p2 PropagateGenerate_WO_0/XOR_WO_1/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1156 PropagateGenerate_WO_0/XOR_WO_1/a_63_n51# PropagateGenerate_WO_0/XOR_WO_1/a_59_n30# gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1157 p2 PropagateGenerate_WO_0/XOR_WO_1/a_51_n59# PropagateGenerate_WO_0/XOR_WO_1/a_63_n51# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1158 PropagateGenerate_WO_0/XOR_WO_1/a_79_n51# a2 p2 Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1159 gnd b2 PropagateGenerate_WO_0/XOR_WO_1/a_79_n51# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1160 PropagateGenerate_WO_0/XOR_WO_0/a_59_n30# b1 PropagateGenerate_WO_0/XOR_WO_0/2INV_1/a_6_87# PropagateGenerate_WO_0/XOR_WO_0/2INV_1/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1161 PropagateGenerate_WO_0/XOR_WO_0/a_59_n30# b1 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1162 PropagateGenerate_WO_0/XOR_WO_0/a_51_n59# a1 vdd PropagateGenerate_WO_0/XOR_WO_0/2INV_0/w_0_81# pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1163 PropagateGenerate_WO_0/XOR_WO_0/a_51_n59# a1 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1164 vdd PropagateGenerate_WO_0/XOR_WO_0/a_51_n59# PropagateGenerate_WO_0/XOR_WO_0/a_56_27# PropagateGenerate_WO_0/XOR_WO_0/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=400 ps=180
M1165 PropagateGenerate_WO_0/XOR_WO_0/a_71_27# PropagateGenerate_WO_0/XOR_WO_0/a_59_n30# vdd PropagateGenerate_WO_0/XOR_WO_0/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1166 p1 a1 PropagateGenerate_WO_0/XOR_WO_0/a_71_27# PropagateGenerate_WO_0/XOR_WO_0/w_50_21# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1167 PropagateGenerate_WO_0/XOR_WO_0/a_56_27# b1 p1 PropagateGenerate_WO_0/XOR_WO_0/w_50_21# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1168 PropagateGenerate_WO_0/XOR_WO_0/a_63_n51# PropagateGenerate_WO_0/XOR_WO_0/a_59_n30# gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1169 p1 PropagateGenerate_WO_0/XOR_WO_0/a_51_n59# PropagateGenerate_WO_0/XOR_WO_0/a_63_n51# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1170 PropagateGenerate_WO_0/XOR_WO_0/a_79_n51# a1 p1 Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1171 gnd b1 PropagateGenerate_WO_0/XOR_WO_0/a_79_n51# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1172 g2_bar a2 vdd PropagateGenerate_WO_0/2AND_WO_1/w_0_0# pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1173 vdd b2 g2_bar PropagateGenerate_WO_0/2AND_WO_1/w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1174 PropagateGenerate_WO_0/2AND_WO_1/a_13_n43# a2 gnd Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1175 g2_bar b2 PropagateGenerate_WO_0/2AND_WO_1/a_13_n43# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1176 g4_bar a4 vdd PropagateGenerate_WO_0/2AND_WO_3/w_0_0# pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1177 vdd b4 g4_bar PropagateGenerate_WO_0/2AND_WO_3/w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1178 PropagateGenerate_WO_0/2AND_WO_3/a_13_n43# a4 gnd Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1179 g4_bar b4 PropagateGenerate_WO_0/2AND_WO_3/a_13_n43# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1180 g1_bar a1 vdd PropagateGenerate_WO_0/2AND_WO_0/w_0_0# pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1181 vdd b1 g1_bar PropagateGenerate_WO_0/2AND_WO_0/w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1182 PropagateGenerate_WO_0/2AND_WO_0/a_13_n43# a1 gnd Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1183 g1_bar b1 PropagateGenerate_WO_0/2AND_WO_0/a_13_n43# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1184 g3_bar a3 vdd PropagateGenerate_WO_0/2AND_WO_2/w_0_0# pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1185 vdd b3 g3_bar PropagateGenerate_WO_0/2AND_WO_2/w_0_0# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1186 PropagateGenerate_WO_0/2AND_WO_2/a_13_n43# a3 gnd Gnd nfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1187 g3_bar b3 PropagateGenerate_WO_0/2AND_WO_2/a_13_n43# Gnd nfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
C0 g4 g3 2.0fF
C1 a3 b3 7.5fF
C2 p2 g2 2.5fF
C3 p2 p3 4.7fF
C4 p2 PropagateGenerate_WO_0/XOR_WO_1/a_56_27# 1.1fF
C5 Carry_WO_0/m1_409_n82# Carry_WO_0/m1_402_n83# 2.3fF
C6 g4 p4 2.0fF
C7 Carry_WO_0/m1_226_n94# g3 1.1fF
C8 g2 p3 6.4fF
C9 g2 Carry_WO_0/m1_63_n31# 1.2fF
C10 SUM_WO_0/XOR_WO_0/a_56_27# s1 1.1fF
C11 g3 p3 2.1fF
C12 c3 p4 2.0fF
C13 p2 g1 10.3fF
C14 a3 b2 2.4fF
C15 a4 b4 12.7fF
C16 a4 b3 5.2fF
C17 vdd g1_bar 1.2fF
C18 PropagateGenerate_WO_0/XOR_WO_3/a_56_27# p4 1.1fF
C19 SUM_WO_0/XOR_WO_3/a_56_27# s4 1.1fF
C20 a1 b1 3.5fF
C21 vdd p3 1.1fF
C22 g3 p4 2.9fF
C23 SUM_WO_0/XOR_WO_2/a_56_27# s3 1.1fF
C24 p4 p3 4.3fF
C25 Carry_WO_0/m1_402_n83# Carry_WO_0/m1_395_n85# 1.5fF
C26 a2 b2 4.8fF
C27 c2 p3 2.0fF
C28 g4 Carry_WO_0/m1_409_n82# 2.9fF
C29 PropagateGenerate_WO_0/XOR_WO_0/a_56_27# p1 1.1fF
C30 gnd p1 2.3fF
C31 PropagateGenerate_WO_0/XOR_WO_2/a_56_27# p3 1.1fF
C32 g1 vdd 1.3fF
C33 SUM_WO_0/XOR_WO_1/a_56_27# s2 1.1fF
C34 g3_bar gnd! 1.8fF
C35 b3 gnd! 5.9fF
C36 PropagateGenerate_WO_0/2AND_WO_2/w_0_0# gnd! 1.0fF
C37 g1_bar gnd! 1.1fF
C38 b1 gnd! 4.1fF
C39 PropagateGenerate_WO_0/2AND_WO_0/w_0_0# gnd! 1.0fF
C40 b4 gnd! 7.4fF
C41 PropagateGenerate_WO_0/2AND_WO_3/w_0_0# gnd! 1.0fF
C42 b2 gnd! 5.8fF
C43 PropagateGenerate_WO_0/2AND_WO_1/w_0_0# gnd! 1.0fF
C44 p1 gnd! 21.1fF
C45 PropagateGenerate_WO_0/XOR_WO_0/w_50_21# gnd! 2.7fF
C46 PropagateGenerate_WO_0/XOR_WO_0/a_51_n59# gnd! 1.6fF
C47 a1 gnd! 3.5fF
C48 PropagateGenerate_WO_0/XOR_WO_1/w_50_21# gnd! 2.7fF
C49 PropagateGenerate_WO_0/XOR_WO_1/a_51_n59# gnd! 1.6fF
C50 a2 gnd! 3.8fF
C51 p3 gnd! 27.0fF
C52 PropagateGenerate_WO_0/XOR_WO_2/w_50_21# gnd! 2.7fF
C53 PropagateGenerate_WO_0/XOR_WO_2/a_51_n59# gnd! 1.6fF
C54 a3 gnd! 4.9fF
C55 p4 gnd! 26.0fF
C56 PropagateGenerate_WO_0/XOR_WO_3/w_50_21# gnd! 2.7fF
C57 PropagateGenerate_WO_0/XOR_WO_3/a_51_n59# gnd! 1.6fF
C58 a4 gnd! 6.5fF
C59 g2_bar gnd! 2.1fF
C60 Carry_WO_0/w_7_77# gnd! 1.0fF
C61 Carry_WO_0/w_38_n91# gnd! 1.8fF
C62 Carry_WO_0/2NAND_WO_1/w_0_0# gnd! 1.0fF
C63 Carry_WO_0/m1_174_23# gnd! 1.2fF
C64 Carry_WO_0/3NAND_WO_0/w_0_0# gnd! 1.3fF
C65 g3 gnd! 15.0fF
C66 Carry_WO_0/2NAND_WO_2/w_0_0# gnd! 1.0fF
C67 Carry_WO_0/m1_395_n85# gnd! 1.5fF
C68 g2 gnd! 16.9fF
C69 Carry_WO_0/3NAND_WO_1/w_0_0# gnd! 1.3fF
C70 vdd gnd! 58.4fF
C71 Carry_WO_0/m1_402_n83# gnd! 1.9fF
C72 Carry_WO_0/3NOR_WO_0/w_1_n3# gnd! 3.1fF
C73 g1 gnd! 19.4fF
C74 p2 gnd! 26.6fF
C75 Carry_WO_0/4NAND_WO_0/w_0_0# gnd! 1.7fF
C76 gnd gnd! 59.6fF
C77 Carry_WO_0/m1_409_n82# gnd! 4.6fF
C78 g4 gnd! 16.3fF
C79 Carry_WO_0/4NOR_WO_0/w_0_0# gnd! 4.6fF
C80 c4 gnd! 5.0fF
C81 s1 gnd! 1.5fF
C82 SUM_WO_0/XOR_WO_0/w_50_21# gnd! 2.7fF
C83 SUM_WO_0/XOR_WO_0/a_51_n59# gnd! 1.6fF
C84 s2 gnd! 1.5fF
C85 SUM_WO_0/XOR_WO_1/w_50_21# gnd! 2.7fF
C86 SUM_WO_0/XOR_WO_1/a_51_n59# gnd! 1.6fF
C87 s3 gnd! 1.5fF
C88 SUM_WO_0/XOR_WO_2/w_50_21# gnd! 2.7fF
C89 SUM_WO_0/XOR_WO_2/a_51_n59# gnd! 1.6fF
C90 c2 gnd! 7.5fF
C91 s4 gnd! 1.6fF
C92 SUM_WO_0/XOR_WO_3/w_50_21# gnd! 2.7fF
C93 SUM_WO_0/XOR_WO_3/a_51_n59# gnd! 1.6fF
C94 c3 gnd! 7.3fF
