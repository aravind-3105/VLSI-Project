* SPICE3 file created from 3AND.ext - technology: scmos
.option scale=0.09u
.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.global gnd vdd

Vdd	vdd	gnd	'SUPPLY'
vdA     A     0 pulse 1.8 0 0ns 100ps 100ps 5ns  30ns
vdB     B     0 pulse 1.8 0 0ns 100ps 100ps 10ns  30ns
vdC     C     0 pulse 1.8 0 0ns 100ps 100ps 20ns  40ns
vd4     D     0 pulse 1.8 0 0ns 100ps 100ps 30ns  50ns

M1000 out D vdd w_0_0# CMOSP w=20 l=2
+  ad=240 pd=104 as=320 ps=152
M1001 vdd C out w_0_0# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 out B vdd w_0_0# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 vdd A out w_0_0# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 a_13_n78# D gnd gnd CMOSN w=40 l=2
+  ad=240 pd=92 as=200 ps=90
M1005 a_21_n78# C a_13_n78# gnd CMOSN w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1006 a_29_n78# B a_21_n78# gnd CMOSN w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1007 out A a_29_n78# gnd CMOSN w=40 l=2
+  ad=280 pd=94 as=0 ps=0
C0 w_0_0# gnd 1.9fF




.tran 1n 80n
.control
set hcopypscolor = 1
set color0=white
set color1=black

run
plot v(A)
plot v(B)
plot v(C)
plot v(D)
plot v(out)
set curplottitle= "Aravind Narayanan-2019102014"
.endc