magic
tech scmos
timestamp 1619561402
<< nwell >>
rect -2 12 126 64
<< ntransistor >>
rect 9 -39 11 -19
rect 45 -39 47 -19
rect 61 -39 63 -19
rect 79 -39 81 -19
rect 91 -39 93 -19
rect 111 -39 113 -19
<< ptransistor >>
rect 11 18 13 58
rect 17 18 19 58
rect 45 18 47 58
rect 81 18 83 58
rect 111 18 113 58
<< ndiffusion >>
rect 6 -39 9 -19
rect 11 -39 30 -19
rect 42 -39 45 -19
rect 47 -39 61 -19
rect 63 -39 66 -19
rect 78 -39 79 -19
rect 81 -39 91 -19
rect 93 -39 96 -19
rect 108 -39 111 -19
rect 113 -39 116 -19
<< pdiffusion >>
rect 8 18 11 58
rect 13 18 17 58
rect 19 18 30 58
rect 42 18 45 58
rect 47 18 58 58
rect 78 18 81 58
rect 83 18 96 58
rect 108 18 111 58
rect 113 18 116 58
<< ndcontact >>
rect 2 -39 6 -19
rect 30 -39 34 -19
rect 38 -39 42 -19
rect 66 -39 70 -19
rect 74 -39 78 -19
rect 96 -39 100 -19
rect 104 -39 108 -19
rect 116 -39 120 -19
<< pdcontact >>
rect 4 18 8 58
rect 30 18 34 58
rect 38 18 42 58
rect 58 18 62 58
rect 74 18 78 58
rect 96 18 100 58
rect 104 18 108 58
rect 116 18 120 58
<< polysilicon >>
rect 11 58 13 61
rect 17 58 19 61
rect 45 58 47 61
rect 81 58 83 61
rect 111 58 113 61
rect 11 9 13 18
rect 11 -5 13 5
rect 9 -7 13 -5
rect 9 -19 11 -7
rect 17 -11 19 18
rect 45 7 47 18
rect 81 9 83 18
rect 111 9 113 18
rect 45 -19 47 3
rect 81 -5 83 5
rect 79 -7 83 -5
rect 61 -19 63 -11
rect 79 -19 81 -7
rect 91 -19 93 -15
rect 111 -19 113 5
rect 9 -42 11 -39
rect 45 -42 47 -39
rect 61 -42 63 -39
rect 79 -42 81 -39
rect 91 -42 93 -39
rect 111 -42 113 -39
<< polycontact >>
rect 9 5 13 9
rect 43 3 47 7
rect 79 5 83 9
rect 109 5 113 9
rect 15 -15 19 -11
rect 59 -11 63 -7
rect 89 -15 93 -11
<< metal1 >>
rect -2 67 126 71
rect 4 58 8 67
rect 38 58 42 67
rect 74 58 78 67
rect 104 58 108 67
rect -2 5 9 9
rect 30 -7 34 18
rect 58 9 62 18
rect 96 9 100 18
rect 116 9 120 18
rect 42 3 43 7
rect 47 3 48 7
rect 58 5 79 9
rect 96 5 109 9
rect 116 5 126 9
rect -2 -15 15 -11
rect 19 -15 22 -11
rect 30 -11 59 -7
rect 30 -19 34 -11
rect 66 -19 70 5
rect 87 -15 89 -11
rect 96 -19 100 5
rect 116 -19 120 5
rect 2 -45 6 -39
rect 38 -45 42 -39
rect 74 -45 78 -39
rect 104 -45 108 -39
rect -2 -49 126 -45
<< m2contact >>
rect 37 3 42 8
rect 48 3 53 8
rect 22 -15 27 -10
rect 82 -15 87 -10
<< metal2 >>
rect 53 3 77 7
rect 37 -11 41 3
rect 27 -15 41 -11
rect 73 -11 77 3
rect 73 -15 82 -11
<< labels >>
rlabel metal1 1 7 1 7 3 D
rlabel metal1 67 -47 67 -47 1 gnd
rlabel metal1 68 69 68 69 5 vdd
rlabel pdiffusion 85 36 85 36 1 g
rlabel metal1 100 7 100 7 1 Q_bar
rlabel metal1 123 7 123 7 7 Q
rlabel metal1 1 -13 1 -13 3 Clk
rlabel pdiffusion 15 38 15 38 1 lp1
rlabel ndiffusion 54 -29 54 -29 1 pn1
rlabel pdiffusion 85 36 85 36 1 lp2
rlabel ndiffusion 85 -29 85 -29 1 pn2
<< end >>
